netcdf census_bmks_lscaled_allyears_1pft_v2bci_201015 {
dimensions:
	datechars = 10 ;
	cens = 5 ;
	confidence = 3 ;
	dclass = 10 ;
variables:
	char census_comp_date(cens, datechars) ;
		census_comp_date:units = "YYYY-MM-DD" ;
	double confidence(confidence) ;
		confidence:units = "-" ;
		confidence:long_name = "Confidence Limit (0.5 is central tendency)" ;
	double dclass(dclass) ;
		dclass:units = "cm" ;
		dclass:long_name = "diameter class lower bound" ;
	float growth_increment_by_size_census(cens, dclass, confidence) ;
		growth_increment_by_size_census:units = "cm yr-1" ;
		growth_increment_by_size_census:_FillValue = -9.e+30f ;
	float mortality_rate_by_size_census(cens, dclass, confidence) ;
		mortality_rate_by_size_census:units = "yr-1" ;
		mortality_rate_by_size_census:_FillValue = -9.e+30f ;
	float basal_area_by_size_census(cens, dclass, confidence) ;
		basal_area_by_size_census:units = "m2 ha-1" ;
		basal_area_by_size_census:_FillValue = -9.e+30f ;
	float abund_by_size_census(cens, dclass, confidence) ;
		abund_by_size_census:units = "ha-1" ;
		abund_by_size_census:_FillValue = -9.e+30f ;
	float new_recruits_by_census(cens, confidence) ;
		new_recruits_by_census:units = "ha-1 yr-1" ;
		new_recruits_by_census:_FillValue = -9.e+30f ;
data:

 census_comp_date =
  "1992-12-04",
  "1996-02-15",
  "2001-03-31",
  "2006-01-24",
  "2011-03-28" ;

 confidence = 0.05, 0.5, 0.95 ;

 dclass = 1, 5, 10, 15, 20, 30, 40, 50, 60, 70 ;

 growth_increment_by_size_census =
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.04445816, 0.04478455, 0.04519255,
  0.1186268, 0.1209223, 0.1233135,
  0.199272, 0.2045639, 0.2100072,
  0.2736962, 0.2849725, 0.2970615,
  0.3608268, 0.3724912, 0.3877899,
  0.459718, 0.4912252, 0.5233973,
  0.5234792, 0.5655937, 0.6066858,
  0.56297, 0.6366103, 0.7059501,
  0.621272, 0.724416, 0.82559,
  0.5205033, 0.6157928, 0.7105577,
  0.05088533, 0.05121573, 0.05147933,
  0.109399, 0.1108382, 0.1126059,
  0.1847841, 0.1904414, 0.1960681,
  0.2634111, 0.2737416, 0.2850287,
  0.3580257, 0.3726051, 0.3912784,
  0.4669248, 0.4971591, 0.5220631,
  0.5683931, 0.6132123, 0.6567709,
  0.6319278, 0.6988293, 0.7700592,
  0.7051731, 0.8064589, 0.8894764,
  0.6098523, 0.6944896, 0.7645153,
  0.05023928, 0.05059886, 0.05093277,
  0.1196327, 0.1214286, 0.1232315,
  0.1903101, 0.1946847, 0.1989897,
  0.268745, 0.2787329, 0.2893034,
  0.3312868, 0.342459, 0.35816,
  0.4460424, 0.475696, 0.5039008,
  0.5961972, 0.6382633, 0.676658,
  0.6422342, 0.730309, 0.8181563,
  0.6522403, 0.7519516, 0.8433989,
  0.4700375, 0.551747, 0.6276686,
  0.06685624, 0.06735875, 0.06792446,
  0.1419129, 0.1443782, 0.1464964,
  0.2103414, 0.2158863, 0.2245796,
  0.2807574, 0.2951189, 0.3087321,
  0.3277684, 0.3384273, 0.3551815,
  0.3921826, 0.4100923, 0.4386931,
  0.5934164, 0.6360927, 0.695725,
  0.6715973, 0.7553835, 0.8426232,
  0.4956519, 0.6228625, 0.7393577,
  0.6600087, 0.749074, 0.8585736 ;

 mortality_rate_by_size_census =
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.0327137, 0.03314307, 0.03357656,
  0.02239591, 0.02327514, 0.02417956,
  0.01981523, 0.02131985, 0.022907,
  0.02014753, 0.02242032, 0.02487598,
  0.01703702, 0.01917311, 0.02149993,
  0.01671729, 0.01984276, 0.02337617,
  0.01691617, 0.02131647, 0.02649747,
  0.0168524, 0.02252323, 0.02946574,
  0.01629143, 0.0237113, 0.03330749,
  0.01141348, 0.01592031, 0.02159974,
  0.03481038, 0.0352572, 0.0357082,
  0.02641532, 0.02735195, 0.02831277,
  0.02303606, 0.02461553, 0.02627316,
  0.02268141, 0.02505292, 0.02760126,
  0.0193477, 0.02157127, 0.02397697,
  0.01787942, 0.02100589, 0.02451489,
  0.01623504, 0.02042744, 0.02535871,
  0.01273592, 0.01761767, 0.02373383,
  0.01167847, 0.01775217, 0.02583284,
  0.01426749, 0.01912284, 0.02508031,
  0.02942921, 0.02985673, 0.03028878,
  0.02445619, 0.02536716, 0.02630284,
  0.02539238, 0.02705725, 0.02880082,
  0.02205013, 0.02444532, 0.02702584,
  0.02099354, 0.0232999, 0.02578684,
  0.0207532, 0.02408113, 0.02778313,
  0.02669517, 0.031864, 0.03772295,
  0.0208854, 0.02698168, 0.0342737,
  0.01678219, 0.02364067, 0.03232554,
  0.01470938, 0.01954513, 0.02544413,
  0.02988691, 0.03032475, 0.03076728,
  0.02229265, 0.02317147, 0.02407557,
  0.02308237, 0.02469914, 0.02639761,
  0.0210059, 0.02337243, 0.02592885,
  0.02213404, 0.02455897, 0.02717311,
  0.0218033, 0.02525922, 0.02909903,
  0.02289226, 0.0277983, 0.03342715,
  0.0163013, 0.02178725, 0.02850311,
  0.01501912, 0.02172543, 0.0303659,
  0.01412233, 0.01887174, 0.02468785 ;

 basal_area_by_size_census =
  1.931018, 1.940975, 1.950133,
  2.225405, 2.248779, 2.273879,
  1.92219, 1.962262, 2.002296,
  1.715394, 1.76141, 1.807169,
  3.267979, 3.357468, 3.45901,
  3.045132, 3.159648, 3.300606,
  2.637784, 2.807464, 2.924115,
  2.470433, 2.624361, 2.817636,
  2.019882, 2.189565, 2.36371,
  9.526007, 10.5451, 11.53241,
  1.80871, 1.816273, 1.824262,
  2.202429, 2.223725, 2.247401,
  1.960385, 1.994427, 2.031735,
  1.716666, 1.769315, 1.816837,
  3.298128, 3.411286, 3.499864,
  3.103253, 3.23317, 3.364491,
  2.737195, 2.868264, 3.008611,
  2.413351, 2.585808, 2.749278,
  2.018413, 2.216191, 2.419536,
  9.61136, 10.50493, 11.31821,
  1.737299, 1.745746, 1.754282,
  2.137507, 2.156969, 2.17911,
  1.942062, 1.97514, 2.009232,
  1.62077, 1.665916, 1.733234,
  3.265824, 3.368378, 3.478692,
  3.127507, 3.257321, 3.362963,
  2.848514, 3.01354, 3.158968,
  2.444252, 2.620933, 2.836995,
  2.164295, 2.380292, 2.598921,
  9.784106, 10.75512, 11.85611,
  1.69751, 1.706401, 1.712822,
  2.13142, 2.153425, 2.176849,
  1.915915, 1.951751, 1.9913,
  1.613146, 1.652208, 1.696462,
  3.222487, 3.292775, 3.387954,
  3.128518, 3.254597, 3.399593,
  2.79244, 2.924162, 3.070788,
  2.452556, 2.629978, 2.783764,
  2.119122, 2.336006, 2.49411,
  9.939273, 10.79014, 11.84353,
  1.730186, 1.737992, 1.747299,
  2.161933, 2.181249, 2.201345,
  1.896171, 1.933703, 1.962673,
  1.645517, 1.690261, 1.728424,
  3.182407, 3.273998, 3.353548,
  3.012088, 3.143782, 3.324067,
  2.655864, 2.816501, 2.968422,
  2.419683, 2.64753, 2.797603,
  2.103261, 2.274916, 2.460685,
  9.959313, 11.04125, 11.7581 ;

 abund_by_size_census =
  4537.82, 4553.52, 4569.22,
  583.8, 589.44, 595.1,
  167.46, 170.5, 173.54,
  73.8, 75.82, 77.86,
  69.66, 71.62, 73.6,
  32.5, 33.84, 35.2,
  16.92, 17.9, 18.88,
  10.52, 11.3, 12.08,
  6.1, 6.7, 7.3,
  11.38, 12.18, 13,
  4145.92, 4160.92, 4175.94,
  581.46, 587.1, 592.74,
  170.68, 173.74, 176.82,
  73.62, 75.64, 77.66,
  70.46, 72.44, 74.42,
  33.04, 34.4, 35.76,
  17.34, 18.32, 19.32,
  10.26, 11.02, 11.8,
  6.2, 6.8, 7.42,
  11.44, 12.24, 13.06,
  3823.4, 3837.78, 3852.22,
  564.18, 569.72, 575.28,
  168.36, 171.4, 174.46,
  69.42, 71.38, 73.36,
  69.98, 71.94, 73.92,
  33.44, 34.8, 36.18,
  18.3, 19.32, 20.34,
  10.4, 11.18, 11.96,
  6.66, 7.28, 7.92,
  11.48, 12.28, 13.1,
  3742.06, 3756.3, 3770.58,
  564.44, 569.98, 575.54,
  165.5, 168.52, 171.54,
  69, 70.96, 72.92,
  68.52, 70.46, 72.42,
  33.3, 34.66, 36.04,
  17.6, 18.6, 19.6,
  10.34, 11.1, 11.88,
  6.44, 7.06, 7.68,
  11.6, 12.42, 13.24,
  3764.64, 3778.92, 3793.24,
  574.36, 579.96, 585.56,
  164.92, 167.92, 170.94,
  71.12, 73.1, 75.1,
  68.16, 70.1, 72.06,
  32.06, 33.4, 34.74,
  16.86, 17.84, 18.82,
  10.4, 11.18, 11.96,
  6.34, 6.94, 7.56,
  12.08, 12.9, 13.74 ;

 new_recruits_by_census =
  _, _, _,
  365.2953, 367.3357, 369.3761,
  308.4773, 310.3102, 312.147,
  326.1532, 328.03, 329.9067,
  346.6721, 348.6211, 350.5701 ;
}
