netcdf BONA_datm {
dimensions:
	time = 365 ;
variables:
	double time(time) ;
		time:units = "days since 2018-01-01 00:00:00.0 -0:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
	double temp_degC(time) ;
		temp_degC:units = "deg_C" ;
		temp_degC:_FillValue = 1.e+32 ;
		temp_degC:long_name = "mean air temperature" ;
	double wind(time) ;
		wind:units = "m/s" ;
		wind:_FillValue = 1.e+32 ;
		wind:long_name = "mean wind speed" ;
	double RH(time) ;
		RH:units = "%" ;
		RH:_FillValue = 1.e+32 ;
		RH:long_name = "mean relative humidity" ;
	double precip(time) ;
		precip:units = "mm" ;
		precip:_FillValue = 1.e+32 ;
		precip:long_name = "mean precipitation" ;
data:

 time = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 
    108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 
    122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 
    136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 
    150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 
    164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 
    178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 
    192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 
    206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 
    220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 
    234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 
    248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 
    262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 
    276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 
    290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 
    304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 
    318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 
    332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 
    346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 
    360, 361, 362, 363, 364, 365 ;

 temp_degC = -15.8853625, -8.00424791666667, -6.54171875, -13.1669997301918, 
    -14.5702412917059, -10.66796875, -16.56529375, -18.2111708333333, 
    -16.0845520833333, -23.4475895833333, -21.16805, -23.7617229166667, 
    -20.3642958333333, -5.87803958333333, -4.14696458333334, 
    -5.79359583333333, 1.17892083333333, -4.71088440547582, 
    -8.48830995010491, -13.908372994484, -24.3034690172092, 
    -25.7048541666667, -22.67045, -31.0578480681818, -30.66270625, 
    -31.385625, -22.3359958333333, -25.8265729166667, -30.3238770833333, 
    -26.8090916666667, -18.7416833333333, -23.8240520833333, 
    -26.5117291666667, -20.0009333333333, -22.28421875, -24.187825, 
    -11.599925, -19.8320791666667, -24.7780625, -20.5686125, 
    -19.5733583333333, -17.8421375, -8.13892291666667, -4.1654125, 
    -5.15173541666666, -4.48501458333334, -7.7082875, -12.2540875, 
    -8.87018541666667, -6.12251458333333, -3.46273125, -5.55024375, 
    -4.4850125, -5.8432875, -16.8338, -15.0979458333333, -14.7962291666667, 
    -12.7161291666667, -17.8616145833333, -24.1731125, -17.8029125, 
    -11.985293586612, -10.0347645833333, -13.5615395833333, -7.40269375, 
    -7.81850833333333, -11.2112270833333, -4.07534166666667, -7.7585875, 
    -8.50188333333333, -5.6252375, -5.12515416666667, -0.843052083333331, 
    -4.27875833333333, -8.28398333333334, -4.562825, -3.15870416666666, 
    -2.15227083333334, -5.11760416666667, -8.29275624999999, -13.94569375, 
    -8.1788875, -6.38291875, -6.91672083333333, -7.36427916666667, 
    -8.74304791666667, -5.37349791666667, -2.89690833333334, 
    -4.17843958333333, -8.75698958333334, -3.09820208333333, -8.6424125, 
    -10.9660770833333, -9.6572625, -4.78563125, -2.70029166666666, 
    -3.55501041666667, -1.20481666666666, -1.42611458333333, 
    1.53700416666667, 4.39426666666667, 2.86008125, 2.65774070518457, 
    -3.32191666666667, -5.26679375, -1.7135375, -0.720177083333328, 
    1.21635625, -1.05647291666667, -4.47515208333333, -6.18699583333333, 
    -2.59409583333333, 2.78564375, 5.90520625, 5.67934375, 3.5104375, 
    2.97360161741553, 2.05670833333334, 3.84908333333333, 2.63283958333333, 
    1.64656875, -0.0187854166666668, 0.817104166666669, 3.84595625000001, 
    6.55111041666666, 3.90850208333333, 3.93313541666667, 6.46284166666667, 
    9.41569791666666, 12.8263020833333, 11.087, 5.49982291666667, 
    6.77506041666667, 9.67847708333333, 6.9785125, 5.50751041666667, 
    5.69528125, 9.68068333333333, 11.4832354166667, 11.7759270833333, 
    11.6714145833333, 11.8845604166667, 11.3163666666667, 8.56831041666667, 
    8.00595208333333, 9.33647916666666, 10.7766375, 9.56567708333333, 
    11.30574375, 11.4224125, 10.4076104166667, 9.45007083333333, 10.80498125, 
    13.6866145833333, 14.5199083333333, 14.7238979166667, 13.6323979166667, 
    14.0971895833333, 12.8116625, 12.8749416666667, 10.4681020833333, 5.9185, 
    6.40264375, 7.14656666666667, 12.22834375, 8.26439791666667, 10.404975, 
    13.1956041666667, 13.7435625, 16.0895083333333, 14.7395645833333, 
    19.9323916666667, 16.56388125, 13.757675, 13.83385, 15.0415833333333, 
    16.9027916666667, 13.8760875, 12.8418729166667, 13.4274145833333, 
    14.1001604166667, 14.7184104166667, 14.0823458333333, 16.37233125, 
    17.0173645833333, 16.5245145833333, 15.9664979166667, 15.5273916666667, 
    18.160525, 14.00126875, 15.6023599431818, 12.7728416666667, 
    10.4698685217101, 10.4559949758477, 12.4248732781991, 15.0491578541393, 
    14.4028174696015, 14.4530131435655, 14.2150691447583, 16.7386256890025, 
    16.7239699482945, 17.01393125, 17.2503030113636, 17.2971063888889, 
    17.228312906586, 17.7055580208333, 17.695549375, 17.3326229166667, 
    14.2576854166667, 15.8327729166667, 18.1488729166667, 19.6728, 
    17.4931145833333, 14.2042395833333, 14.38230625, 14.7370375, 
    13.6791541666667, 12.89563125, 11.5731020833333, 9.95230833333333, 
    8.97619375, 10.1454791666667, 9.5207875, 13.6811666666667, 
    13.6827895833333, 11.6422354166667, 10.2341916666667, 9.61988668499711, 
    10.0983791666667, 10.18543125, 10.2075145833333, 14.3359979166667, 
    14.500875, 10.79938125, 8.82695625, 10.76464375, 10.0734625, 
    7.47197708333334, 11.0637708333333, 9.96030416666666, 9.29078125, 
    6.66794166666666, 5.20359166666667, 3.8382875, 9.17527916666667, 
    9.44221041666667, 8.55998541666667, 9.0582375, 8.8325625, 7.72569375, 
    6.8042125, 3.80459791666667, 4.21940833333333, 7.47067291666666, 
    9.44323680555556, 11.4285434944356, 6.04151750848501, 9.2017, 8.65715, 
    8.48204791666667, 8.68761041666667, 8.96666666666667, 6.887775, 7.503075, 
    6.61481458333334, 6.00895208333333, 6.29355833333333, 7.16717291666666, 
    5.685375, 3.9766, 2.98968333333333, 5.69374791666667, 4.45229583333333, 
    9.8773375, 6.02090416666667, 3.22587291666667, 6.13019583333333, 
    3.65342708333333, 3.60305416666666, 0.695983333333333, -6.90489166666666, 
    -5.66236458333333, 1.44356666666667, 2.06094375, 0.472895833333331, 
    3.17698541666667, 3.16847708333334, 0.0680645833333339, 6.2587125, 
    1.93069791666667, 1.74074472588541, 0.886237499999998, 1.44490625, 
    -0.152743749999999, -0.648883333333329, 3.18370208333333, 
    5.15241666666666, 0.132816666666667, 3.31381352623535, 0.260862347003314, 
    -1.82671458333333, -7.86547291666667, -14.3570875, -17.9095520833333, 
    -12.1169083333333, -12.8819041666667, -13.9185458333333, -17.2963875, 
    -16.9147229166667, -16.9385770833333, -14.6810104166667, -11.59009375, 
    -13.7702134635051, -7.81819375, -7.00809166666666, -3.9286875, 
    -8.33709791666667, -9.7756875, -15.01895, -18.034275, -14.5888708333333, 
    -11.9094020833333, -6.24861458333333, -7.31516458333333, 
    -9.05141401473542, -12.2443035958836, -10.6629854166667, 
    -12.7676291666667, -13.8588458333333, -10.377575, -6.63719791666667, 
    -11.24510625, -10.6075484659408, -11.0599607272988, -14.5099782808519, 
    -6.15478125, -7.04216875, -7.17923541666666, -8.87692708333333, 
    -7.41575416666667, -5.54239637516659, -5.070225, -9.82926458333333, 
    -17.4377208333333, -16.1333541666667, -15.4386375, -19.1745395833333, 
    -22.51086875, -24.0732916666667, -24.4737916666667, -23.8599791666667, 
    -19.2512014785882, -15.9184657592801, -21.6648351113431, 
    -28.0273020833333, -20.6911020833333, -23.1696770833333, -19.50170625, 
    -20.80709375, -25.6126791666667, -20.96830625, -20.2791979166667, 
    -20.2325270833333, -18.01815, -5.371525 ;

 wind = 1.35104498704351, 2.08949516902496, 1.62617868411728, 
    1.16804301843004, 1.2127458440856, 2.46711609113151, 1.91280873172156, 
    2.13626437791593, 4.30180884890822, 1.83456246407361, 0.724973003105274, 
    1.04372658987038, 1.04616640681873, 2.7683820258648, 1.65560189648208, 
    1.5888305222356, 1.5496090387044, 1.02454354893772, 0.753944342170138, 
    0.86979969117542, 1.06667276675782, 0.689670279085623, 0.7015528789836, 
    1.07351848750609, 0.939077198318063, 1.01026196987924, 1.37058665909938, 
    1.22578465643676, 1.02747575696571, 1.25830149805772, 2.92267984610739, 
    2.12497471735855, 1.10348042652042, 2.09000949323901, 1.08579756032526, 
    0.919104938072392, 2.11825824737449, 1.73820410992777, 1.41088343143339, 
    1.27530399307781, 1.45107060332125, 1.02347268579637, 0.897756572396289, 
    2.33661423001597, 1.5020063348565, 1.36220498679989, 1.4493539397013, 
    0.992660541763114, 1.11809182494485, 0.947937513253106, 1.91121110092576, 
    1.65910477834014, 0.847061351531248, 4.72181657964166, 1.87604047700597, 
    3.26751115139342, 1.2414452518488, 3.03095898721745, 1.57638819232172, 
    1.56574374812233, 1.21989561361954, 0.80018646656083, 0.851196505932279, 
    1.32790453188043, 1.01831447717511, 1.66987034581667, 1.82910087128428, 
    2.58474279899724, 1.4435489097042, 1.80591311219037, 1.73167227906065, 
    2.00651245238741, 1.73262623478503, 1.69748938033609, 1.55608821503264, 
    0.693639943069844, 1.20557793340422, 2.03585908104218, 2.3325535140728, 
    1.76916584069615, 1.76017225420306, 2.86887712496725, 2.92038001228639, 
    3.31633998586928, 3.57609842886948, 2.77785016858992, 1.38444767376755, 
    1.35968768638328, 1.57540265968347, 1.97682966694803, 1.72049460280601, 
    2.13702105298261, 3.69196934290738, 5.59635682114149, 4.44596513893986, 
    3.99780375293149, 1.98341805307411, 3.24012237658596, 2.94110458420808, 
    3.72437721424, 2.49984109647243, 1.73288979034058, 2.48880095129735, 
    2.63342061116561, 3.34448970303495, 3.21988403837379, 3.29387271795257, 
    3.42317791743869, 4.33101962788799, 4.18986070582149, 3.10394570181152, 
    2.27128136284336, 2.43267654065479, 2.83578098781156, 2.54500238224905, 
    2.45168643560425, 1.98798715964644, 1.80697634481247, 1.52539497885874, 
    1.81329532298571, 1.74455841653835, 2.76624195406167, 2.0116048106718, 
    2.90532972546352, 2.5505764744865, 2.09875071608883, 2.25924462667128, 
    2.42467970562167, 3.60106880430249, 3.6127469849426, 3.26842752683565, 
    2.27713495912224, 1.8916283479851, 2.60313801413039, 1.83353373592423, 
    2.20002830538862, 2.12175902855918, 2.95191773132701, 3.26005362967998, 
    3.11822666856092, 2.53989711828801, 2.27377305760654, 1.61736259654549, 
    1.77510629265785, 1.71535446639568, 2.30691451763929, 3.7179201931684, 
    2.74045189613215, 2.13864577975239, 2.22500520441643, 1.87598770530102, 
    1.58600994736732, 1.98988307048643, 2.04257016985857, 2.1478664946626, 
    2.95652483294815, 2.72322256528867, 2.36266976447533, 1.92199688016794, 
    2.22622928672235, 2.0553500358375, 2.14872073505129, 1.61421509762019, 
    1.37813667625117, 2.80373904668155, 2.60581264266545, 1.08689087601803, 
    1.52581630497534, 1.89985337181252, 2.15113247538138, 1.49931585109399, 
    1.72067308685215, 1.90659865459096, 2.65887653813281, 2.15729972939868, 
    1.85769271711276, 2.34811394552521, 1.87886118906296, 1.5922486590805, 
    1.54401827607087, 1.95868195974977, 1.48147252629583, 2.27243880361733, 
    3.22106055943792, 3.07812667506569, 2.27851504055495, 2.15224841968031, 
    1.97545753562323, 2.46831682455074, 1.64416021309526, 1.67467397146474, 
    1.81982493248812, 1.97125645521715, 1.98796864958172, 1.93570094901821, 
    1.98597361993952, 1.87051331309195, 1.93518483829357, 2.12865859141426, 
    2.36098988774533, 2.37576657844245, 2.25534350347082, 2.09048739074949, 
    2.09481102005675, 2.11971647925077, 2.03325445402714, 2.04074365774322, 
    1.78165448606055, 1.73892945462948, 1.68271213450255, 1.87851481336595, 
    1.64719736650922, 2.15857993037233, 1.33655331792662, 1.38785098116001, 
    1.33219517090681, 1.83700852787976, 1.58753228890419, 1.6156040401072, 
    1.5393988577831, 2.25063634521709, 1.78678539915238, 1.65472840709951, 
    1.57393529536852, 1.54630766732464, 1.01320466863119, 1.64506966429602, 
    2.29675465266114, 2.09327447974972, 1.69369897489124, 1.73693368323878, 
    1.13534618050603, 0.940469335160978, 2.22859138852265, 1.04102543423641, 
    1.08423100474904, 1.95510120057377, 1.25865540044275, 1.78385678397405, 
    2.51202567442054, 1.95938395930954, 1.86669250450768, 2.09450446388996, 
    1.86562223977151, 3.05509806543078, 2.19616734794738, 2.28455867124734, 
    1.76715218664216, 1.26227462407645, 2.47539214462938, 2.63512378763309, 
    1.55951746511678, 1.47140736474889, 1.52043606249522, 1.80699474828031, 
    1.74649362904518, 2.59205475827751, 1.44586602294259, 1.51362050188372, 
    1.11411603805553, 1.21143009242423, 1.1185160826794, 0.880894330993611, 
    1.01947646945244, 1.18147595443397, 0.916401659715889, 1.86443346769077, 
    1.70314362203642, 1.33597572312888, 2.05040330246927, 3.07765765660415, 
    2.61183917767856, 2.22384362288424, 2.98885643247321, 2.38251103343681, 
    1.74450611968903, 2.87314942792755, 2.08773109609107, 1.15860206425236, 
    2.557547669307, 1.74011894661137, 2.00503978516226, 2.5419954585817, 
    1.26730572256631, 1.25139318335366, 1.87267207420954, 1.06018863206294, 
    2.3059484132581, 2.11576003810471, 1.11408087902195, 1.44060484600806, 
    3.03497174213073, 1.48557091058754, 1.7369594246392, 1.62840563428649, 
    4.43388957077842, 2.31149512115411, 1.77063419980347, 1.95403695842576, 
    0.987482007027187, 1.48129178472961, 1.43760509488812, 1.37730236310328, 
    1.56174668973575, 1.57021582160659, 1.93080005576915, 1.79312010596229, 
    1.07838509885058, 1.36265053335107, 1.44613650263056, 1.19611617115427, 
    0.942185818384539, 1.51246932044015, 0.697346325747528, 1.93008792557045, 
    1.67759670069453, 3.36526983442148, 2.2867640322133, 1.9854045317936, 
    1.18579100072544, 1.11802419288228, 1.00585709687195, 1.15904589665577, 
    1.00960081266109, 1.10370217640821, 0.618418086643147, 0.740663847300886, 
    1.18138316974673, 1.11663927683065, 1.25171692977564, 1.3628126823256, 
    1.1765693768274, 0.830028638892579, 0.930643618506227, 1.45090876368238, 
    1.99374513973832, 1.09687936099784, 1.37254919664542, 1.36926762555664, 
    1.38533816100251, 1.42426876606307, 1.25876888476348, 0.924877687280245, 
    1.63190643917753, 1.25382371515097, 0.942715645094827, 0.828210591532498, 
    1.42234058643138, 0.867099100289516, 0.942715645094828, 
    0.846034491379465, 0.729909083285592, 0.952437772284083, 
    0.994566990104184, 1.12878635713361, 0.87006975026401, 0.891944536439833, 
    2.38213058728166, 1.98352337252223, 1.23221898806374, 0.911658849906932, 
    1.17199581130808, 1.26273566507445, 1.15768267961279, 1.95301377922511 ;

 RH = 83.9229166666667, 90.088125, 90.5679166666667, 86.9397916666667, 
    85.396875, 86.8727083333333, 82.0077083333333, 79.2354166666667, 
    66.940625, 76.1652083333333, 79.1864583333333, 77.363125, 
    79.3447916666667, 83.8402083333333, 93.361875, 92.0877083333333, 
    99.0113882751379, 94.86625, 91.6922916666667, 86.8070833333333, 
    78.6633333333333, 78.0410416666667, 80.5066666666667, 74.5050492424242, 
    74.440625, 73.799375, 80.4227083333333, 76.7477083333333, 
    73.7495833333333, 76.4229166666667, 79.4972916666667, 76.8770833333333, 
    74.9975, 78.9422916666667, 77.6160416666667, 76.5402083333333, 
    82.7191666666667, 78.936875, 75.965, 78.3897916666667, 79.1691666666667, 
    82.6264583333333, 91.2333333333333, 92.3858333333333, 92.9079166666667, 
    92.8270833333333, 89.23125, 87.490625, 89.451875, 91.896875, 
    92.4622916666667, 88.39125, 93.7720833333333, 86.0513182997257, 
    79.453125, 78.5639583333333, 82.6483333333333, 84.23625, 
    83.4622916666667, 72.4345833333333, 77.4495833333333, 85.1766666666667, 
    85.91, 79.8116179930599, 87.7097916666667, 83.19625, 75.54875, 
    71.1466666666667, 82.5625, 79.77125, 77.4275, 78.59, 85.4091666666667, 
    86.92625, 85.84, 89.2589583333333, 88.2597916666667, 93.10125, 
    89.3095833333333, 87.9252083333333, 82.9835416666667, 73.2227083333333, 
    62.3435416666667, 51.6664583333333, 49.6464583333333, 55.0397916666667, 
    61.7845833333333, 74.7516666666667, 75.09875, 72.995, 82.215, 61.741875, 
    57.6272916666667, 51.8535416666667, 48.1447916666667, 52.911875, 
    62.3077083333333, 58.5279166666667, 61.6560416666667, 51.3227083333333, 
    59.7704166666667, 69.1883333333333, 70.9302083333333, 65.3875, 
    56.9216666666667, 45.6522916666667, 53.7454166666667, 48.533125, 
    42.624375, 51.8145833333333, 67.9233333333333, 63.424375, 
    54.8447916666667, 63.4452083333333, 67.2647916666667, 61.6541666666667, 
    67.5870833333333, 63.39375, 67.6133333333333, 91.3295833333333, 
    88.8695833333333, 77.361875, 60.3375, 59.7175, 56.4133333333333, 
    61.681875, 63.0491666666667, 51.358125, 51.0095833333333, 49.278125, 
    59.0779166666667, 71.6535416666667, 55.793125, 48.7020833333333, 
    67.4097916666667, 75.7347916666667, 62.540625, 54.9729166666667, 
    67.34125, 58.1302083333333, 71.7027083333333, 63.0045833333333, 
    74.6208333333333, 89.8775363938355, 85.4758333333333, 68.8008333333333, 
    55.605, 51.2116666666667, 47.2479364920843, 66.20125, 65.38125, 
    85.1052083333333, 66.9708333333333, 56.9808333333333, 59.0889583333333, 
    60.7295833333333, 73.529375, 54.7716666666667, 61.56125, 65.059375, 
    79.8258333333333, 89.5722751206075, 74.15875, 69.041875, 
    61.1754166666667, 55.735, 78.9610416666667, 73.9335416666667, 
    64.4333333333333, 63.86, 62.4145833333333, 53.6475, 81.246867767761, 
    72.1239583333333, 60.1445833333333, 57.5610416666667, 57.778125, 
    77.986875, 82.0408333333333, 82.5760416666667, 79.2566666666667, 
    88.1072916666667, 87.5270833333333, 65.510625, 56.2333333333333, 
    70.0333333333333, 72.03375, 69.7429166666667, 65.7775, 76.4191666666667, 
    58.6040340909091, 81.3285416666667, 97.0545347222222, 97.05034375, 
    84.8332438257658, 71.966571428333, 73.2949953758565, 72.8253323662111, 
    77.1662185236468, 65.43809375, 65.4177465277778, 65.3152083333333, 
    65.0251183712121, 64.9350173611111, 69.2598429659498, 69.6211319444444, 
    69.69375, 71.4316959451015, 86.0589583333333, 69.0595833333333, 
    63.4154166666667, 61.8235416666667, 74.7772916666667, 84.4741666666667, 
    84.0730113636364, 88.25, 95.018801549995, 96.5268390376113, 
    89.8802083333333, 81.8089583333333, 67.4225, 74.509375, 72.9914583333333, 
    75.3047916666667, 79.001875, 95.4531876140769, 96.6060442314667, 
    88.1294253589018, 86.2560416666667, 86.505, 76.9085416666667, 
    79.1545833333333, 89.9033333333333, 81.985625, 85.627253139478, 
    92.4745906511784, 90.0966666666667, 88.196875, 95.5325, 93.1863678795947, 
    87.18125, 91.4520833333333, 94.0778737322737, 89.8364583333333, 
    93.1276753333575, 91.2629166666667, 87.5670833333333, 89.264375, 92.9525, 
    85.308125, 74.1485416666667, 77.350625, 79.0291666666667, 
    76.7135416666667, 82.2736111111111, 80.4329166666667, 68.2945833333333, 
    60.2410416666667, 74.7272916666667, 85.2910416666667, 79.868125, 
    91.9084073880472, 96.2539583333333, 96.3810416666667, 97.715, 
    98.7077932743805, 96.3586448943785, 96.258125, 96.6611226933847, 
    86.1164583333333, 79.0507920063241, 67.2091143009064, 65.8260416666667, 
    57.2285416666667, 56.3670833333333, 68.0833333333333, 58.5127083333333, 
    64.6245833333333, 68.6697916666667, 57.3591666666667, 69.535625, 
    68.6470833333333, 59.286875, 94.9520833333333, 96.4877083333333, 
    97.8737689169178, 95.0422296811714, 89.6875, 91.3411431310437, 97.1875, 
    95.346056470449, 88.8879166666667, 94.8577083333333, 95.9656377076798, 
    92.3810416666667, 80.9870833333333, 84.6033333333333, 91.4122916666667, 
    88.6691666666667, 95.161875, 92.8735416666667, 84.931875, 83.52625, 
    80.9479166666667, 85.1022916666667, 83.71125, 82.8225, 80.29, 80.500625, 
    81.2191666666667, 83.6945833333333, 87.23375, 85.0194952173809, 
    91.1097916666667, 89.5310416666667, 91.2560416666667, 83.8408333333333, 
    80.92375, 80.2527083333333, 80.9052083333333, 83.925625, 
    86.8416666666667, 91.4985416666667, 91.239375, 90.6316666666667, 
    87.1660416666667, 88.3952083333333, 86.1591666666667, 84.8114583333333, 
    87.8802602195128, 89.4320833333333, 84.7183333333333, 89.4635416666667, 
    88.11125, 84.6225, 90.6166666666667, 91.0566666666667, 90.048125, 
    88.8460416666667, 88.8916666666667, 92.22125, 92.84, 89.3458333333333, 
    80.63875, 81.3070833333333, 84.8616666666667, 81.56875, 77.915625, 
    77.9702083333333, 77.1258333333333, 78.3377083333333, 81.9504703952504, 
    83.195, 79.0089583333333, 73.849375, 80.3914583333333, 76.475, 
    78.1110416666667, 77.6539583333333, 75.8645833333333, 79.22375, 
    79.291875, 79.074375, 82.3997916666667, 89.9479166666667 ;

 precip = 0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 1.21286391042609, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.886760629555732, 0.886760629555732, 0.886760629555732, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.825667622993205, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.95638982935677, 0.782319326582488, 0.782319326582488, 1.10777020822857, 
    0.782319326582488, 4.13199120000743, 0.782319326582488, 1.04274776361249, 
    3.67480213630066, 0.869015919403921, 0.956389829356769, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    1.41290157593212, 0.744176026474195, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.842483528867979, 0.6, 0.89, 1.5, 1.13, 0.77, 0.9, 1.34, 0.64, 0.68, 
    1.03, 0.86, 0.91, 1.23, 1.91, 1.04, 0.75, 0.619999999999999, 0.63, 2.04, 
    1.2, 1.21, 0.800000000000001, 2.31, 1.2, 1.05, 1.24, 0.583983781370185, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 1.87814495765951, 
    0.737790167821228, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.889386722093501, 1.13, 
    0.89593512548074, 0.802838318706262, 0.769386722093501, 0.69, 0.4, 
    0.959999999999999, 1.01, 1.23, 1.09, 0.96, 0.67, 0.57, 0.366903193225522, 
    2.12, 4.11, 2.93, 1.17, 0.72, 0.83, 0.31, 0.85, 0.68, 0.7, 5.23, 2.09, 
    0.13, 0.41, 0.82, 1.18, 0.52, 0.74, 0.490000000000001, 1.02, 1.38, 0.58, 
    0.83, 1.93, 0.63, 0.62, 4.33, 1.38, 0.73, 2.35, 0.53, 0.28, 0.63, 1.65, 
    0.67, 1.27, 1.4, 1.01, 0.9, 0.223451596612761, 0.79, 1.4, 1.07, 0.23, 
    0.56, 0.81, 0.540000000000001, 1.15, 3.82, 4.46, 5.3, 1.64, 2, 0.44, 
    1.57, 1.33, 1.18, 1.46, 0.959999999999999, 1.04, 0.5, 1.19, 1.08, 0.48, 
    0.59, 0.87, 0.24, 0.86, 0.42, 0.47, 0.24, 0.47, 0.29, 1.27, 0.6, 0.37, 
    0.81, 0.25, 0.21, 0.51, 0.34, 0.91, 0.570000000000001, 0.43, 0.46, 
    0.0799999999999999, 0.18672579830638, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 0.802838318706262, 
    0.802838318706262, 0.802838318706262, 1.08230613394884, 0.45, 
    0.418144957659511, 0.802838318706262, 0.731773949191413, 0.89, 0.72, 
    0.15, 0.04, 0.66, 0.37, 0.42, 0.11, 0.38, 0.52, 0.94, 0.77, 
    0.44005462120265, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 
    0.782319326582488, 0.782319326582488, 0.782319326582488, 0.782319326582488 ;
}
