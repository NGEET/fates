netcdf param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908 {
dimensions:
	fates_NCWD = 4 ;
	fates_history_age_bins = 7 ;
	fates_history_coage_bins = 2 ;
	fates_history_height_bins = 6 ;
	fates_history_size_bins = 13 ;
	fates_hydr_organs = 4 ;
	fates_leafage_class = 1 ;
	fates_litterclass = 6 ;
	fates_pft = 3 ;
	fates_prt_organs = 6 ;
	fates_string_length = 60 ;
variables:
	double fates_history_sizeclass_bin_edges(fates_history_size_bins) ;
		fates_history_sizeclass_bin_edges:units = "cm" ;
		fates_history_sizeclass_bin_edges:long_name = "Lower edges for DBH size class bins used in size-resolved cohort history output" ;
	double fates_history_ageclass_bin_edges(fates_history_age_bins) ;
		fates_history_ageclass_bin_edges:units = "yr" ;
		fates_history_ageclass_bin_edges:long_name = "Lower edges for age class bins used in age-resolved patch history output" ;
	char fates_prt_organ_name(fates_prt_organs, fates_string_length) ;
		fates_prt_organ_name:units = "unitless - string" ;
		fates_prt_organ_name:long_name = "Plant organ name (order must match PRTGenericMod.F90)" ;
	double fates_prt_alloc_priority(fates_prt_organs, fates_pft) ;
		fates_prt_alloc_priority:units = "index (0-fates_prt_organs)" ;
		fates_prt_alloc_priority:long_name = "Priority order for allocation" ;
	double fates_prt_nitr_stoich_p1(fates_prt_organs, fates_pft) ;
		fates_prt_nitr_stoich_p1:units = "(gN/gC)" ;
		fates_prt_nitr_stoich_p1:long_name = "nitrogen stoichiometry, parameter 1" ;
	double fates_prt_nitr_stoich_p2(fates_prt_organs, fates_pft) ;
		fates_prt_nitr_stoich_p2:units = "(gN/gC)" ;
		fates_prt_nitr_stoich_p2:long_name = "nitrogen stoichiometry, parameter 2" ;
	double fates_prt_phos_stoich_p1(fates_prt_organs, fates_pft) ;
		fates_prt_phos_stoich_p1:units = "(gP/gC)" ;
		fates_prt_phos_stoich_p1:long_name = "phosphorous stoichiometry, parameter 1" ;
	double fates_prt_phos_stoich_p2(fates_prt_organs, fates_pft) ;
		fates_prt_phos_stoich_p2:units = "(gP/gC)" ;
		fates_prt_phos_stoich_p2:long_name = "phosphorous stoichiometry, parameter 2" ;
	double fates_turnover_carb_retrans(fates_prt_organs, fates_pft) ;
		fates_turnover_carb_retrans:units = "-" ;
		fates_turnover_carb_retrans:long_name = "retranslocation fraction of carbon in turnover" ;
	double fates_turnover_nitr_retrans(fates_prt_organs, fates_pft) ;
		fates_turnover_nitr_retrans:units = "-" ;
		fates_turnover_nitr_retrans:long_name = "retranslocation fraction of nitrogen in turnover" ;
	double fates_turnover_phos_retrans(fates_prt_organs, fates_pft) ;
		fates_turnover_phos_retrans:units = "-" ;
		fates_turnover_phos_retrans:long_name = "retranslocation fraction of phosphorous in turnover, parameter 1" ;
	double fates_fire_FBD(fates_litterclass) ;
		fates_fire_FBD:units = "NA" ;
		fates_fire_FBD:long_name = "spitfire parameter related to fuel bulk density, see SFMain.F90" ;
	double fates_fire_SAV(fates_litterclass) ;
		fates_fire_SAV:units = "NA" ;
		fates_fire_SAV:long_name = "spitfire parameter related to surface area to volume ratio, see SFMain.F90" ;
	double fates_fire_low_moisture_Coeff(fates_litterclass) ;
		fates_fire_low_moisture_Coeff:units = "NA" ;
		fates_fire_low_moisture_Coeff:long_name = "spitfire parameter, equation B1 Thonicke et al 2010" ;
	double fates_fire_low_moisture_Slope(fates_litterclass) ;
		fates_fire_low_moisture_Slope:units = "NA" ;
		fates_fire_low_moisture_Slope:long_name = "spitfire parameter, equation B1 Thonicke et al 2010" ;
	double fates_fire_mid_moisture(fates_litterclass) ;
		fates_fire_mid_moisture:units = "NA" ;
		fates_fire_mid_moisture:long_name = "spitfire litter moisture threshold to be considered medium dry" ;
	double fates_fire_mid_moisture_Coeff(fates_litterclass) ;
		fates_fire_mid_moisture_Coeff:units = "NA" ;
		fates_fire_mid_moisture_Coeff:long_name = "spitfire parameter, equation B1 Thonicke et al 2010" ;
	double fates_fire_mid_moisture_Slope(fates_litterclass) ;
		fates_fire_mid_moisture_Slope:units = "NA" ;
		fates_fire_mid_moisture_Slope:long_name = "spitfire parameter, equation B1 Thonicke et al 2010" ;
	double fates_fire_min_moisture(fates_litterclass) ;
		fates_fire_min_moisture:units = "NA" ;
		fates_fire_min_moisture:long_name = "spitfire litter moisture threshold to be considered very dry" ;
	double fates_history_height_bin_edges(fates_history_height_bins) ;
		fates_history_height_bin_edges:units = "m" ;
		fates_history_height_bin_edges:long_name = "Lower edges for height bins used in height-resolved history output" ;
	double fates_max_decomp(fates_litterclass) ;
		fates_max_decomp:units = "yr-1" ;
		fates_max_decomp:long_name = "maximum rate of litter & CWD transfer from non-decomposing class into decomposing class" ;
	double fates_hydr_avuln_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_avuln_node:units = "unitless" ;
		fates_hydr_avuln_node:long_name = "xylem vulnerability curve shape parameter" ;
	double fates_hydr_epsil_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_epsil_node:units = "MPa" ;
		fates_hydr_epsil_node:long_name = "bulk elastic modulus" ;
	double fates_hydr_fcap_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_fcap_node:units = "unitless" ;
		fates_hydr_fcap_node:long_name = "fraction of non-residual water that is capillary in source" ;
	double fates_hydr_kmax_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_kmax_node:units = "kg/MPa/m/s" ;
		fates_hydr_kmax_node:long_name = "maximum xylem conductivity per unit conducting xylem area" ;
	double fates_hydr_p50_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_p50_node:units = "MPa" ;
		fates_hydr_p50_node:long_name = "xylem water potential at 50% loss of conductivity" ;
	double fates_hydr_pinot_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_pinot_node:units = "MPa" ;
		fates_hydr_pinot_node:long_name = "osmotic potential at full turgor" ;
	double fates_hydr_pitlp_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_pitlp_node:units = "MPa" ;
		fates_hydr_pitlp_node:long_name = "turgor loss point" ;
	double fates_hydr_resid_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_resid_node:units = "cm3/cm3" ;
		fates_hydr_resid_node:long_name = "residual water conent" ;
	double fates_hydr_thetas_node(fates_hydr_organs, fates_pft) ;
		fates_hydr_thetas_node:units = "cm3/cm3" ;
		fates_hydr_thetas_node:long_name = "saturated water content" ;
	double fates_CWD_frac(fates_NCWD) ;
		fates_CWD_frac:units = "fraction" ;
		fates_CWD_frac:long_name = "fraction of woody (bdead+bsw) biomass destined for CWD pool" ;
	char fates_pftname(fates_pft, fates_string_length) ;
		fates_pftname:units = "unitless - string" ;
		fates_pftname:long_name = "Description of plant type" ;
	double fates_alloc_storage_cushion(fates_pft) ;
		fates_alloc_storage_cushion:units = "fraction" ;
		fates_alloc_storage_cushion:long_name = "maximum size of storage C pool, relative to maximum size of leaf C pool" ;
	double fates_allom_agb1(fates_pft) ;
		fates_allom_agb1:units = "variable" ;
		fates_allom_agb1:long_name = "Parameter 1 for agb allometry" ;
	double fates_allom_agb2(fates_pft) ;
		fates_allom_agb2:units = "variable" ;
		fates_allom_agb2:long_name = "Parameter 2 for agb allometry" ;
	double fates_allom_agb3(fates_pft) ;
		fates_allom_agb3:units = "variable" ;
		fates_allom_agb3:long_name = "Parameter 3 for agb allometry" ;
	double fates_allom_agb4(fates_pft) ;
		fates_allom_agb4:units = "variable" ;
		fates_allom_agb4:long_name = "Parameter 4 for agb allometry" ;
	double fates_allom_agb_frac(fates_pft) ;
		fates_allom_agb_frac:units = "fraction" ;
		fates_allom_agb_frac:long_name = "Fraction of woody biomass that is above ground" ;
	double fates_allom_amode(fates_pft) ;
		fates_allom_amode:units = "index" ;
		fates_allom_amode:long_name = "AGB allometry function index." ;
	double fates_allom_blca_expnt_diff(fates_pft) ;
		fates_allom_blca_expnt_diff:units = "unitless" ;
		fates_allom_blca_expnt_diff:long_name = "difference between allometric DBH:bleaf and DBH:crown area exponents" ;
	double fates_allom_cmode(fates_pft) ;
		fates_allom_cmode:units = "index" ;
		fates_allom_cmode:long_name = "coarse root biomass allometry function index." ;
	double fates_allom_d2bl1(fates_pft) ;
		fates_allom_d2bl1:units = "variable" ;
		fates_allom_d2bl1:long_name = "Parameter 1 for d2bl allometry" ;
	double fates_allom_d2bl2(fates_pft) ;
		fates_allom_d2bl2:units = "variable" ;
		fates_allom_d2bl2:long_name = "Parameter 2 for d2bl allometry" ;
	double fates_allom_d2bl3(fates_pft) ;
		fates_allom_d2bl3:units = "unitless" ;
		fates_allom_d2bl3:long_name = "Parameter 3 for d2bl allometry" ;
	double fates_allom_d2ca_coefficient_max(fates_pft) ;
		fates_allom_d2ca_coefficient_max:units = "m2 cm^(-1/beta)" ;
		fates_allom_d2ca_coefficient_max:long_name = "max (savanna) dbh to area multiplier factor where: area = n*d2ca_coeff*dbh^beta" ;
	double fates_allom_d2ca_coefficient_min(fates_pft) ;
		fates_allom_d2ca_coefficient_min:units = "m2 cm^(-1/beta)" ;
		fates_allom_d2ca_coefficient_min:long_name = "min (forest) dbh to area multiplier factor where: area = n*d2ca_coeff*dbh^beta" ;
	double fates_allom_d2h1(fates_pft) ;
		fates_allom_d2h1:units = "variable" ;
		fates_allom_d2h1:long_name = "Parameter 1 for d2h allometry (intercept, or c)" ;
	double fates_allom_d2h2(fates_pft) ;
		fates_allom_d2h2:units = "variable" ;
		fates_allom_d2h2:long_name = "Parameter 2 for d2h allometry (slope, or m)" ;
	double fates_allom_d2h3(fates_pft) ;
		fates_allom_d2h3:units = "variable" ;
		fates_allom_d2h3:long_name = "Parameter 3 for d2h allometry (optional)" ;
	double fates_allom_dbh_maxheight(fates_pft) ;
		fates_allom_dbh_maxheight:units = "cm" ;
		fates_allom_dbh_maxheight:long_name = "the diameter (if any) corresponding to maximum height, diameters may increase beyond this" ;
	double fates_allom_fmode(fates_pft) ;
		fates_allom_fmode:units = "index" ;
		fates_allom_fmode:long_name = "fine root biomass allometry function index." ;
	double fates_allom_frbstor_repro(fates_pft) ;
		fates_allom_frbstor_repro:units = "fraction" ;
		fates_allom_frbstor_repro:long_name = "fraction of bstore goes to reproduction after plant dies" ;
	double fates_allom_hmode(fates_pft) ;
		fates_allom_hmode:units = "index" ;
		fates_allom_hmode:long_name = "height allometry function index." ;
	double fates_allom_l2fr(fates_pft) ;
		fates_allom_l2fr:units = "gC/gC" ;
		fates_allom_l2fr:long_name = "Allocation parameter: fine root C per leaf C" ;
	double fates_allom_la_per_sa_int(fates_pft) ;
		fates_allom_la_per_sa_int:units = "m2/cm2" ;
		fates_allom_la_per_sa_int:long_name = "Leaf area per sapwood area, intercept" ;
	double fates_allom_la_per_sa_slp(fates_pft) ;
		fates_allom_la_per_sa_slp:units = "m2/cm2/m" ;
		fates_allom_la_per_sa_slp:long_name = "Leaf area per sapwood area rate of change with height, slope (optional)" ;
	double fates_allom_lmode(fates_pft) ;
		fates_allom_lmode:units = "index" ;
		fates_allom_lmode:long_name = "leaf biomass allometry function index." ;
	double fates_allom_sai_scaler(fates_pft) ;
		fates_allom_sai_scaler:units = "m2/m2" ;
		fates_allom_sai_scaler:long_name = "allometric ratio of SAI per LAI" ;
	double fates_allom_smode(fates_pft) ;
		fates_allom_smode:units = "index" ;
		fates_allom_smode:long_name = "sapwood allometry function index." ;
	double fates_allom_stmode(fates_pft) ;
		fates_allom_stmode:units = "index" ;
		fates_allom_stmode:long_name = "storage allometry function index." ;
	double fates_branch_turnover(fates_pft) ;
		fates_branch_turnover:units = "yr" ;
		fates_branch_turnover:long_name = "turnover time of branches" ;
	double fates_c2b(fates_pft) ;
		fates_c2b:units = "ratio" ;
		fates_c2b:long_name = "Carbon to biomass multiplier of bulk structural tissues" ;
	double fates_displar(fates_pft) ;
		fates_displar:units = "unitless" ;
		fates_displar:long_name = "Ratio of displacement height to canopy top height" ;
	double fates_eca_alpha_ptase(fates_pft) ;
		fates_eca_alpha_ptase:units = "g/m3" ;
		fates_eca_alpha_ptase:long_name = "fraction of P from ptase activity sent directly to plant (ECA)" ;
	double fates_eca_decompmicc(fates_pft) ;
		fates_eca_decompmicc:units = "gC/m3" ;
		fates_eca_decompmicc:long_name = "mean soil microbial decomposer biomass (ECA)" ;
	double fates_eca_km_nh4(fates_pft) ;
		fates_eca_km_nh4:units = "gN/m3" ;
		fates_eca_km_nh4:long_name = "half-saturation constant for plant nh4 uptake (ECA)" ;
	double fates_eca_km_no3(fates_pft) ;
		fates_eca_km_no3:units = "gN/m3" ;
		fates_eca_km_no3:long_name = "half-saturation constant for plant no3 uptake (ECA)" ;
	double fates_eca_km_p(fates_pft) ;
		fates_eca_km_p:units = "gP/m3" ;
		fates_eca_km_p:long_name = "half-saturation constant for plant p uptake (ECA)" ;
	double fates_eca_km_ptase(fates_pft) ;
		fates_eca_km_ptase:units = "gP/m3" ;
		fates_eca_km_ptase:long_name = "half-saturation constant for biochemical P (ECA)" ;
	double fates_eca_lambda_ptase(fates_pft) ;
		fates_eca_lambda_ptase:units = "g/m3" ;
		fates_eca_lambda_ptase:long_name = "critical value for biochemical production (ECA)" ;
	double fates_eca_vmax_nh4(fates_pft) ;
		fates_eca_vmax_nh4:units = "gN/gC/s" ;
		fates_eca_vmax_nh4:long_name = "maximum production rate for plant nh4 uptake (ECA)" ;
	double fates_eca_vmax_no3(fates_pft) ;
		fates_eca_vmax_no3:units = "gN/gC/s" ;
		fates_eca_vmax_no3:long_name = "maximum production rate for plant no3 uptake (ECA)" ;
	double fates_eca_vmax_p(fates_pft) ;
		fates_eca_vmax_p:units = "gP/gC/s" ;
		fates_eca_vmax_p:long_name = "maximum production rate for plant p uptake (ECA)" ;
	double fates_eca_vmax_ptase(fates_pft) ;
		fates_eca_vmax_ptase:units = "gP/m2/s" ;
		fates_eca_vmax_ptase:long_name = "maximum production rate for biochemical P (per m2) (ECA)" ;
	double fates_fire_alpha_SH(fates_pft) ;
		fates_fire_alpha_SH:units = "NA" ;
		fates_fire_alpha_SH:long_name = "spitfire parameter, alpha scorch height, Equation 16 Thonicke et al 2010" ;
	double fates_fire_bark_scaler(fates_pft) ;
		fates_fire_bark_scaler:units = "fraction" ;
		fates_fire_bark_scaler:long_name = "the thickness of a cohorts bark as a fraction of its dbh" ;
	double fates_fire_crown_depth_frac(fates_pft) ;
		fates_fire_crown_depth_frac:units = "fraction" ;
		fates_fire_crown_depth_frac:long_name = "the depth of a cohorts crown as a fraction of its height" ;
	double fates_fire_crown_kill(fates_pft) ;
		fates_fire_crown_kill:units = "NA" ;
		fates_fire_crown_kill:long_name = "fire parameter, see equation 22 in Thonicke et al 2010" ;
	double fates_fnrt_prof_a(fates_pft) ;
		fates_fnrt_prof_a:units = "unitless" ;
		fates_fnrt_prof_a:long_name = "Fine root profile function, parameter a" ;
	double fates_fnrt_prof_b(fates_pft) ;
		fates_fnrt_prof_b:units = "unitless" ;
		fates_fnrt_prof_b:long_name = "Fine root profile function, parameter b" ;
	double fates_fnrt_prof_mode(fates_pft) ;
		fates_fnrt_prof_mode:units = "index" ;
		fates_fnrt_prof_mode:long_name = "Index to select fine root profile function: 1) Jackson Beta, 2) 1-param exponential 3) 2-param exponential" ;
	double fates_fr_fcel(fates_pft) ;
		fates_fr_fcel:units = "fraction" ;
		fates_fr_fcel:long_name = "Fine root litter cellulose fraction" ;
	double fates_fr_flab(fates_pft) ;
		fates_fr_flab:units = "fraction" ;
		fates_fr_flab:long_name = "Fine root litter labile fraction" ;
	double fates_fr_flig(fates_pft) ;
		fates_fr_flig:units = "fraction" ;
		fates_fr_flig:long_name = "Fine root litter lignin fraction" ;
	double fates_grperc(fates_pft) ;
		fates_grperc:units = "unitless" ;
		fates_grperc:long_name = "Growth respiration factor" ;
	double fates_hydr_avuln_gs(fates_pft) ;
		fates_hydr_avuln_gs:units = "unitless" ;
		fates_hydr_avuln_gs:long_name = "shape parameter for stomatal control of water vapor exiting leaf" ;
	double fates_hydr_p50_gs(fates_pft) ;
		fates_hydr_p50_gs:units = "MPa" ;
		fates_hydr_p50_gs:long_name = "water potential at 50% loss of stomatal conductance" ;
	double fates_hydr_p_taper(fates_pft) ;
		fates_hydr_p_taper:units = "unitless" ;
		fates_hydr_p_taper:long_name = "xylem taper exponent" ;
	double fates_hydr_rfrac_stem(fates_pft) ;
		fates_hydr_rfrac_stem:units = "fraction" ;
		fates_hydr_rfrac_stem:long_name = "fraction of total tree resistance from troot to canopy" ;
	double fates_hydr_rs2(fates_pft) ;
		fates_hydr_rs2:units = "m" ;
		fates_hydr_rs2:long_name = "absorbing root radius" ;
	double fates_hydr_srl(fates_pft) ;
		fates_hydr_srl:units = "m g-1" ;
		fates_hydr_srl:long_name = "specific root length" ;
	double fates_leaf_c3psn(fates_pft) ;
		fates_leaf_c3psn:units = "flag" ;
		fates_leaf_c3psn:long_name = "Photosynthetic pathway (1=c3, 0=c4)" ;
	double fates_leaf_clumping_index(fates_pft) ;
		fates_leaf_clumping_index:units = "fraction (0-1)" ;
		fates_leaf_clumping_index:long_name = "factor describing how much self-occlusion of leaf scattering elements decreases light interception" ;
	double fates_leaf_diameter(fates_pft) ;
		fates_leaf_diameter:units = "m" ;
		fates_leaf_diameter:long_name = "Characteristic leaf dimension" ;
	double fates_leaf_jmaxha(fates_pft) ;
		fates_leaf_jmaxha:units = "J/mol" ;
		fates_leaf_jmaxha:long_name = "activation energy for jmax" ;
	double fates_leaf_jmaxhd(fates_pft) ;
		fates_leaf_jmaxhd:units = "J/mol" ;
		fates_leaf_jmaxhd:long_name = "deactivation energy for jmax" ;
	double fates_leaf_jmaxse(fates_pft) ;
		fates_leaf_jmaxse:units = "J/mol/K" ;
		fates_leaf_jmaxse:long_name = "entropy term for jmax" ;
	double fates_leaf_slamax(fates_pft) ;
		fates_leaf_slamax:units = "m^2/gC" ;
		fates_leaf_slamax:long_name = "Maximum Specific Leaf Area (SLA), even if under a dense canopy" ;
	double fates_leaf_slatop(fates_pft) ;
		fates_leaf_slatop:units = "m^2/gC" ;
		fates_leaf_slatop:long_name = "Specific Leaf Area (SLA) at top of canopy, projected area basis" ;
	double fates_leaf_stomatal_intercept(fates_pft) ;
		fates_leaf_stomatal_intercept:units = "umol H2O/m**2/s" ;
		fates_leaf_stomatal_intercept:long_name = "Minimum unstressed stomatal conductance for Ball-Berry model and Medlyn model" ;
	double fates_leaf_stomatal_slope_ballberry(fates_pft) ;
		fates_leaf_stomatal_slope_ballberry:units = "unitless" ;
		fates_leaf_stomatal_slope_ballberry:long_name = "stomatal slope parameter, as per Ball-Berry" ;
	double fates_leaf_stomatal_slope_medlyn(fates_pft) ;
		fates_leaf_stomatal_slope_medlyn:units = "KPa**0.5" ;
		fates_leaf_stomatal_slope_medlyn:long_name = "stomatal slope parameter, as per Medlyn" ;
	double fates_leaf_stor_priority(fates_pft) ;
		fates_leaf_stor_priority:units = "unitless" ;
		fates_leaf_stor_priority:long_name = "factor governing priority of replacing storage with NPP" ;
	double fates_leaf_tpuha(fates_pft) ;
		fates_leaf_tpuha:units = "J/mol" ;
		fates_leaf_tpuha:long_name = "activation energy for tpu" ;
	double fates_leaf_tpuhd(fates_pft) ;
		fates_leaf_tpuhd:units = "J/mol" ;
		fates_leaf_tpuhd:long_name = "deactivation energy for tpu" ;
	double fates_leaf_tpuse(fates_pft) ;
		fates_leaf_tpuse:units = "J/mol/K" ;
		fates_leaf_tpuse:long_name = "entropy term for tpu" ;
	double fates_leaf_vcmaxha(fates_pft) ;
		fates_leaf_vcmaxha:units = "J/mol" ;
		fates_leaf_vcmaxha:long_name = "activation energy for vcmax" ;
	double fates_leaf_vcmaxhd(fates_pft) ;
		fates_leaf_vcmaxhd:units = "J/mol" ;
		fates_leaf_vcmaxhd:long_name = "deactivation energy for vcmax" ;
	double fates_leaf_vcmaxse(fates_pft) ;
		fates_leaf_vcmaxse:units = "J/mol/K" ;
		fates_leaf_vcmaxse:long_name = "entropy term for vcmax" ;
	double fates_leaf_xl(fates_pft) ;
		fates_leaf_xl:units = "unitless" ;
		fates_leaf_xl:long_name = "Leaf/stem orientation index" ;
	double fates_lf_fcel(fates_pft) ;
		fates_lf_fcel:units = "fraction" ;
		fates_lf_fcel:long_name = "Leaf litter cellulose fraction" ;
	double fates_lf_flab(fates_pft) ;
		fates_lf_flab:units = "fraction" ;
		fates_lf_flab:long_name = "Leaf litter labile fraction" ;
	double fates_lf_flig(fates_pft) ;
		fates_lf_flig:units = "fraction" ;
		fates_lf_flig:long_name = "Leaf litter lignin fraction" ;
	double fates_maintresp_reduction_curvature(fates_pft) ;
		fates_maintresp_reduction_curvature:units = "unitless (0-1)" ;
		fates_maintresp_reduction_curvature:long_name = "curvature of MR reduction as f(carbon storage), 1=linear, 0=very curved" ;
	double fates_maintresp_reduction_intercept(fates_pft) ;
		fates_maintresp_reduction_intercept:units = "unitless (0-1)" ;
		fates_maintresp_reduction_intercept:long_name = "intercept of MR reduction as f(carbon storage), 0=no throttling, 1=max throttling" ;
	double fates_mort_bmort(fates_pft) ;
		fates_mort_bmort:units = "1/yr" ;
		fates_mort_bmort:long_name = "background mortality rate" ;
	double fates_mort_freezetol(fates_pft) ;
		fates_mort_freezetol:units = "degrees C" ;
		fates_mort_freezetol:long_name = "minimum temperature tolerance" ;
	double fates_mort_hf_flc_threshold(fates_pft) ;
		fates_mort_hf_flc_threshold:units = "fraction" ;
		fates_mort_hf_flc_threshold:long_name = "plant fractional loss of conductivity at which drought mortality begins for hydraulic model" ;
	double fates_mort_hf_sm_threshold(fates_pft) ;
		fates_mort_hf_sm_threshold:units = "unitless" ;
		fates_mort_hf_sm_threshold:long_name = "soil moisture (btran units) at which drought mortality begins for non-hydraulic model" ;
	double fates_mort_ip_age_senescence(fates_pft) ;
		fates_mort_ip_age_senescence:units = "years" ;
		fates_mort_ip_age_senescence:long_name = "Mortality cohort age senescence inflection point. If _ this mortality term is off. Setting this value turns on age dependent mortality. " ;
	double fates_mort_ip_size_senescence(fates_pft) ;
		fates_mort_ip_size_senescence:units = "dbh cm" ;
		fates_mort_ip_size_senescence:long_name = "Mortality dbh senescence inflection point. If _ this mortality term is off. Setting this value turns on size dependent mortality" ;
	double fates_mort_r_age_senescence(fates_pft) ;
		fates_mort_r_age_senescence:units = "mortality rate year^-1" ;
		fates_mort_r_age_senescence:long_name = "Mortality age senescence rate of change. Sensible range is around 0.03-0.06. Larger values givesteeper mortality curves." ;
	double fates_mort_r_size_senescence(fates_pft) ;
		fates_mort_r_size_senescence:units = "mortality rate dbh^-1" ;
		fates_mort_r_size_senescence:long_name = "Mortality dbh senescence rate of change. Sensible range is around 0.03-0.06. Larger values give steeper mortality curves." ;
	double fates_mort_scalar_coldstress(fates_pft) ;
		fates_mort_scalar_coldstress:units = "1/yr" ;
		fates_mort_scalar_coldstress:long_name = "maximum mortality rate from cold stress" ;
	double fates_mort_scalar_cstarvation(fates_pft) ;
		fates_mort_scalar_cstarvation:units = "1/yr" ;
		fates_mort_scalar_cstarvation:long_name = "maximum mortality rate from carbon starvation" ;
	double fates_mort_scalar_hydrfailure(fates_pft) ;
		fates_mort_scalar_hydrfailure:units = "1/yr" ;
		fates_mort_scalar_hydrfailure:long_name = "maximum mortality rate from hydraulic failure" ;
	double fates_nfix1(fates_pft) ;
		fates_nfix1:units = "NA" ;
		fates_nfix1:long_name = "place-holder for future n-fixation parameter (NOT IMPLEMENTED)" ;
	double fates_nfix2(fates_pft) ;
		fates_nfix2:units = "NA" ;
		fates_nfix2:long_name = "place-holder for future n-fixation parameter (NOT IMPLEMENTED)" ;
	double fates_phen_cold_size_threshold(fates_pft) ;
		fates_phen_cold_size_threshold:units = "cm" ;
		fates_phen_cold_size_threshold:long_name = "the dbh size above which will lead to phenology-related stem and leaf drop" ;
	double fates_phen_evergreen(fates_pft) ;
		fates_phen_evergreen:units = "logical flag" ;
		fates_phen_evergreen:long_name = "Binary flag for evergreen leaf habit" ;
	double fates_phen_season_decid(fates_pft) ;
		fates_phen_season_decid:units = "logical flag" ;
		fates_phen_season_decid:long_name = "Binary flag for seasonal-deciduous leaf habit" ;
	double fates_phen_stem_drop_fraction(fates_pft) ;
		fates_phen_stem_drop_fraction:units = "fraction" ;
		fates_phen_stem_drop_fraction:long_name = "fraction of stems to drop for non-woody species during drought/cold" ;
	double fates_phen_stress_decid(fates_pft) ;
		fates_phen_stress_decid:units = "logical flag" ;
		fates_phen_stress_decid:long_name = "Binary flag for stress-deciduous leaf habit" ;
	double fates_phenflush_fraction(fates_pft) ;
		fates_phenflush_fraction:units = "fraction" ;
		fates_phenflush_fraction:long_name = "Upon bud-burst, the maximum fraction of storage carbon used for flushing leaves" ;
	double fates_prescribed_mortality_canopy(fates_pft) ;
		fates_prescribed_mortality_canopy:units = "1/yr" ;
		fates_prescribed_mortality_canopy:long_name = "mortality rate of canopy trees for prescribed physiology mode" ;
	double fates_prescribed_mortality_understory(fates_pft) ;
		fates_prescribed_mortality_understory:units = "1/yr" ;
		fates_prescribed_mortality_understory:long_name = "mortality rate of understory trees for prescribed physiology mode" ;
	double fates_prescribed_npp_canopy(fates_pft) ;
		fates_prescribed_npp_canopy:units = "kgC / m^2 / yr" ;
		fates_prescribed_npp_canopy:long_name = "NPP per unit crown area of canopy trees for prescribed physiology mode" ;
	double fates_prescribed_npp_understory(fates_pft) ;
		fates_prescribed_npp_understory:units = "kgC / m^2 / yr" ;
		fates_prescribed_npp_understory:long_name = "NPP per unit crown area of understory trees for prescribed physiology mode" ;
	double fates_prescribed_nuptake(fates_pft) ;
		fates_prescribed_nuptake:units = "fraction" ;
		fates_prescribed_nuptake:long_name = "Nitrogen uptake flux as fraction of NPP demand. 0=fully coupled simulation" ;
	double fates_prescribed_puptake(fates_pft) ;
		fates_prescribed_puptake:units = "fraction" ;
		fates_prescribed_puptake:long_name = "Phosphorus uptake flux as fraction of NPP demand. 0=fully coupled simulation" ;
	double fates_prescribed_recruitment(fates_pft) ;
		fates_prescribed_recruitment:units = "n/yr" ;
		fates_prescribed_recruitment:long_name = "recruitment rate for prescribed physiology mode" ;
	double fates_recruit_hgt_min(fates_pft) ;
		fates_recruit_hgt_min:units = "m" ;
		fates_recruit_hgt_min:long_name = "the minimum height (ie starting height) of a newly recruited plant" ;
	double fates_recruit_initd(fates_pft) ;
		fates_recruit_initd:units = "stems/m2" ;
		fates_recruit_initd:long_name = "initial seedling density for a cold-start near-bare-ground simulation" ;
	double fates_rholnir(fates_pft) ;
		fates_rholnir:units = "fraction" ;
		fates_rholnir:long_name = "Leaf reflectance: near-IR" ;
	double fates_rholvis(fates_pft) ;
		fates_rholvis:units = "fraction" ;
		fates_rholvis:long_name = "Leaf reflectance: visible" ;
	double fates_rhosnir(fates_pft) ;
		fates_rhosnir:units = "fraction" ;
		fates_rhosnir:long_name = "Stem reflectance: near-IR" ;
	double fates_rhosvis(fates_pft) ;
		fates_rhosvis:units = "fraction" ;
		fates_rhosvis:long_name = "Stem reflectance: visible" ;
	double fates_root_long(fates_pft) ;
		fates_root_long:units = "yr" ;
		fates_root_long:long_name = "root longevity (alternatively, turnover time)" ;
	double fates_seed_alloc(fates_pft) ;
		fates_seed_alloc:units = "fraction" ;
		fates_seed_alloc:long_name = "fraction of available carbon balance allocated to seeds" ;
	double fates_seed_alloc_mature(fates_pft) ;
		fates_seed_alloc_mature:units = "fraction" ;
		fates_seed_alloc_mature:long_name = "fraction of available carbon balance allocated to seeds in mature plants (adds to fates_seed_alloc)" ;
	double fates_seed_dbh_repro_threshold(fates_pft) ;
		fates_seed_dbh_repro_threshold:units = "cm" ;
		fates_seed_dbh_repro_threshold:long_name = "the diameter (if any) where the plant will start extra clonal allocation to the seed pool" ;
	double fates_seed_decay_rate(fates_pft) ;
		fates_seed_decay_rate:units = "yr-1" ;
		fates_seed_decay_rate:long_name = "fraction of seeds that decay per year" ;
	double fates_seed_germination_rate(fates_pft) ;
		fates_seed_germination_rate:units = "yr-1" ;
		fates_seed_germination_rate:long_name = "fraction of seeds that germinate per year" ;
	double fates_seed_suppl(fates_pft) ;
		fates_seed_suppl:units = "KgC/m2/yr" ;
		fates_seed_suppl:long_name = "Supplemental external seed rain source term (non-mass conserving)" ;
	double fates_senleaf_long_fdrought(fates_pft) ;
		fates_senleaf_long_fdrought:units = "unitless[0-1]" ;
		fates_senleaf_long_fdrought:long_name = "multiplication factor for leaf longevity of senescent leaves during drought" ;
	double fates_smpsc(fates_pft) ;
		fates_smpsc:units = "mm" ;
		fates_smpsc:long_name = "Soil water potential at full stomatal closure" ;
	double fates_smpso(fates_pft) ;
		fates_smpso:units = "mm" ;
		fates_smpso:long_name = "Soil water potential at full stomatal opening" ;
	double fates_taulnir(fates_pft) ;
		fates_taulnir:units = "fraction" ;
		fates_taulnir:long_name = "Leaf transmittance: near-IR" ;
	double fates_taulvis(fates_pft) ;
		fates_taulvis:units = "fraction" ;
		fates_taulvis:long_name = "Leaf transmittance: visible" ;
	double fates_tausnir(fates_pft) ;
		fates_tausnir:units = "fraction" ;
		fates_tausnir:long_name = "Stem transmittance: near-IR" ;
	double fates_tausvis(fates_pft) ;
		fates_tausvis:units = "fraction" ;
		fates_tausvis:long_name = "Stem transmittance: visible" ;
	double fates_trim_inc(fates_pft) ;
		fates_trim_inc:units = "m2/m2" ;
		fates_trim_inc:long_name = "Arbitrary incremental change in trimming function." ;
	double fates_trim_limit(fates_pft) ;
		fates_trim_limit:units = "m2/m2" ;
		fates_trim_limit:long_name = "Arbitrary limit to reductions in leaf area with stress" ;
	double fates_turnover_retrans_mode(fates_pft) ;
		fates_turnover_retrans_mode:units = "index" ;
		fates_turnover_retrans_mode:long_name = "retranslocation method for leaf/fineroot turnover." ;
	double fates_wood_density(fates_pft) ;
		fates_wood_density:units = "g/cm3" ;
		fates_wood_density:long_name = "mean density of woody tissue in plant" ;
	double fates_woody(fates_pft) ;
		fates_woody:units = "logical flag" ;
		fates_woody:long_name = "Binary woody lifeform flag" ;
	double fates_z0mr(fates_pft) ;
		fates_z0mr:units = "unitless" ;
		fates_z0mr:long_name = "Ratio of momentum roughness length to canopy top height" ;
	double fates_history_coageclass_bin_edges(fates_history_coage_bins) ;
		fates_history_coageclass_bin_edges:units = "years" ;
		fates_history_coageclass_bin_edges:long_name = "Lower edges for cohort age class bins used in cohort age resolved history output" ;
	double fates_leaf_long(fates_leafage_class, fates_pft) ;
		fates_leaf_long:units = "yr" ;
		fates_leaf_long:long_name = "Leaf longevity (ie turnover timescale)" ;
	double fates_leaf_vcmax25top(fates_leafage_class, fates_pft) ;
		fates_leaf_vcmax25top:units = "umol CO2/m^2/s" ;
		fates_leaf_vcmax25top:long_name = "maximum carboxylation rate of Rub. at 25C, canopy top" ;
	double fates_base_mr_20 ;
		fates_base_mr_20:units = "gC/gN/s" ;
		fates_base_mr_20:long_name = "Base maintenance respiration rate for plant tissues, using Ryan 1991" ;
	double fates_canopy_closure_thresh ;
		fates_canopy_closure_thresh:units = "unitless" ;
		fates_canopy_closure_thresh:long_name = "tree canopy coverage at which crown area allometry changes from savanna to forest value" ;
	double fates_cohort_age_fusion_tol ;
		fates_cohort_age_fusion_tol:units = "unitless" ;
		fates_cohort_age_fusion_tol:long_name = "minimum fraction in differece in cohort age between cohorts." ;
	double fates_cohort_size_fusion_tol ;
		fates_cohort_size_fusion_tol:units = "unitless" ;
		fates_cohort_size_fusion_tol:long_name = "minimum fraction in difference in dbh between cohorts" ;
	double fates_comp_excln ;
		fates_comp_excln:units = "none" ;
		fates_comp_excln:long_name = "IF POSITIVE: weighting factor (exponent on dbh) for canopy layer exclusion and promotion, IF NEGATIVE: switch to use deterministic height sorting" ;
	double fates_cwd_fcel ;
		fates_cwd_fcel:units = "unitless" ;
		fates_cwd_fcel:long_name = "Cellulose fraction for CWD" ;
	double fates_cwd_flig ;
		fates_cwd_flig:units = "unitless" ;
		fates_cwd_flig:long_name = "Lignin fraction of coarse woody debris" ;
	double fates_eca_plant_escalar ;
		fates_eca_plant_escalar:units = "" ;
		fates_eca_plant_escalar:long_name = "scaling factor for plant fine root biomass to calculate nutrient carrier enzyme abundance (ECA)" ;
	double fates_fire_active_crown_fire ;
		fates_fire_active_crown_fire:units = "0 or 1" ;
		fates_fire_active_crown_fire:long_name = "flag, 1=active crown fire 0=no active crown fire" ;
	double fates_fire_cg_strikes ;
		fates_fire_cg_strikes:units = "fraction (0-1)" ;
		fates_fire_cg_strikes:long_name = "fraction of cloud to ground lightning strikes" ;
	double fates_fire_drying_ratio ;
		fates_fire_drying_ratio:units = "NA" ;
		fates_fire_drying_ratio:long_name = "spitfire parameter, fire drying ratio for fuel moisture, alpha_FMC EQ 6 Thonicke et al 2010" ;
	double fates_fire_durat_slope ;
		fates_fire_durat_slope:units = "NA" ;
		fates_fire_durat_slope:long_name = "spitfire parameter, fire max duration slope, Equation 14 Thonicke et al 2010" ;
	double fates_fire_fdi_a ;
		fates_fire_fdi_a:units = "NA" ;
		fates_fire_fdi_a:long_name = "spitfire parameter, fire danger index,  EQ 5 Thonicke et al 2010" ;
	double fates_fire_fdi_alpha ;
		fates_fire_fdi_alpha:units = "NA" ;
		fates_fire_fdi_alpha:long_name = "spitfire parameter, EQ 7 Venevsky et al. GCB 2002,(modified EQ 8 Thonicke et al. 2010) " ;
	double fates_fire_fdi_b ;
		fates_fire_fdi_b:units = "NA" ;
		fates_fire_fdi_b:long_name = "spitfire parameter, fire danger index, EQ 5 Thonicke et al 2010 " ;
	double fates_fire_fuel_energy ;
		fates_fire_fuel_energy:units = "kJ/kg" ;
		fates_fire_fuel_energy:long_name = "spitfire parameter, heat content of fuel" ;
	double fates_fire_max_durat ;
		fates_fire_max_durat:units = "minutes" ;
		fates_fire_max_durat:long_name = "spitfire parameter, fire maximum duration, Equation 14 Thonicke et al 2010" ;
	double fates_fire_miner_damp ;
		fates_fire_miner_damp:units = "NA" ;
		fates_fire_miner_damp:long_name = "spitfire parameter, mineral-dampening coefficient EQ A1 Thonicke et al 2010 " ;
	double fates_fire_miner_total ;
		fates_fire_miner_total:units = "fraction" ;
		fates_fire_miner_total:long_name = "spitfire parameter, total mineral content, Table A1 Thonicke et al 2010" ;
	double fates_fire_nignitions ;
		fates_fire_nignitions:units = "ignitions per year per km2" ;
		fates_fire_nignitions:long_name = "number of annual ignitions per square km" ;
	double fates_fire_part_dens ;
		fates_fire_part_dens:units = "kg/m2" ;
		fates_fire_part_dens:long_name = "spitfire parameter, oven dry particle density, Table A1 Thonicke et al 2010" ;
	double fates_fire_threshold ;
		fates_fire_threshold:units = "kW/m" ;
		fates_fire_threshold:long_name = "spitfire parameter, fire intensity threshold for tracking fires that spread" ;
	double fates_hydr_kmax_rsurf1 ;
		fates_hydr_kmax_rsurf1:units = "kg water/m2 root area/Mpa/s" ;
		fates_hydr_kmax_rsurf1:long_name = "maximum conducitivity for unit root surface (into root)" ;
	double fates_hydr_kmax_rsurf2 ;
		fates_hydr_kmax_rsurf2:units = "kg water/m2 root area/Mpa/s" ;
		fates_hydr_kmax_rsurf2:long_name = "maximum conducitivity for unit root surface (out of root)" ;
	double fates_hydr_psi0 ;
		fates_hydr_psi0:units = "MPa" ;
		fates_hydr_psi0:long_name = "sapwood water potential at saturation" ;
	double fates_hydr_psicap ;
		fates_hydr_psicap:units = "MPa" ;
		fates_hydr_psicap:long_name = "sapwood water potential at which capillary reserves exhausted" ;
	double fates_init_litter ;
		fates_init_litter:units = "NA" ;
		fates_init_litter:long_name = "Initialization value for litter pool in cold-start (NOT USED)" ;
	double fates_leaf_stomatal_model ;
		fates_leaf_stomatal_model:units = "unitless" ;
		fates_leaf_stomatal_model:long_name = "switch for choosing between Ball-Berry (1) stomatal conductance model and Medlyn (2) model" ;
	double fates_logging_coll_under_frac ;
		fates_logging_coll_under_frac:units = "fraction" ;
		fates_logging_coll_under_frac:long_name = "Fraction of stems killed in the understory when logging generates disturbance" ;
	double fates_logging_collateral_frac ;
		fates_logging_collateral_frac:units = "fraction" ;
		fates_logging_collateral_frac:long_name = "Fraction of large stems in upperstory that die from logging collateral damage" ;
	double fates_logging_dbhmax ;
		fates_logging_dbhmax:units = "cm" ;
		fates_logging_dbhmax:long_name = "Maximum dbh below which logging is applied (unset values flag this to be unused)" ;
	double fates_logging_dbhmax_infra ;
		fates_logging_dbhmax_infra:units = "cm" ;
		fates_logging_dbhmax_infra:long_name = "Tree diameter, above which infrastructure from logging does not impact damage or mortality." ;
	double fates_logging_dbhmin ;
		fates_logging_dbhmin:units = "cm" ;
		fates_logging_dbhmin:long_name = "Minimum dbh at which logging is applied" ;
	double fates_logging_direct_frac ;
		fates_logging_direct_frac:units = "fraction" ;
		fates_logging_direct_frac:long_name = "Fraction of stems logged directly per event" ;
	double fates_logging_event_code ;
		fates_logging_event_code:units = "unitless" ;
		fates_logging_event_code:long_name = "Integer code that options how logging events are structured" ;
	double fates_logging_export_frac ;
		fates_logging_export_frac:units = "fraction" ;
		fates_logging_export_frac:long_name = "fraction of trunk product being shipped offsite, the leftovers will be left onsite as large CWD" ;
	double fates_logging_mechanical_frac ;
		fates_logging_mechanical_frac:units = "fraction" ;
		fates_logging_mechanical_frac:long_name = "Fraction of stems killed due infrastructure an other mechanical means" ;
	double fates_mort_disturb_frac ;
		fates_mort_disturb_frac:units = "fraction" ;
		fates_mort_disturb_frac:long_name = "fraction of canopy mortality that results in disturbance (i.e. transfer of area from new to old patch)" ;
	double fates_mort_understorey_death ;
		fates_mort_understorey_death:units = "fraction" ;
		fates_mort_understorey_death:long_name = "fraction of plants in understorey cohort impacted by overstorey tree-fall" ;
	double fates_patch_fusion_tol ;
		fates_patch_fusion_tol:units = "unitless" ;
		fates_patch_fusion_tol:long_name = "minimum fraction in difference in profiles between patches" ;
	double fates_phen_a ;
		fates_phen_a:units = "none" ;
		fates_phen_a:long_name = "GDD accumulation function, intercept parameter: gdd_thesh = a + b exp(c*ncd)" ;
	double fates_phen_b ;
		fates_phen_b:units = "none" ;
		fates_phen_b:long_name = "GDD accumulation function, multiplier parameter: gdd_thesh = a + b exp(c*ncd)" ;
	double fates_phen_c ;
		fates_phen_c:units = "none" ;
		fates_phen_c:long_name = "GDD accumulation function, exponent parameter: gdd_thesh = a + b exp(c*ncd)" ;
	double fates_phen_chiltemp ;
		fates_phen_chiltemp:units = "degrees C" ;
		fates_phen_chiltemp:long_name = "chilling day counting threshold for vegetation" ;
	double fates_phen_coldtemp ;
		fates_phen_coldtemp:units = "degrees C" ;
		fates_phen_coldtemp:long_name = "vegetation temperature exceedance that flags a cold-day for leaf-drop" ;
	double fates_phen_doff_time ;
		fates_phen_doff_time:units = "days" ;
		fates_phen_doff_time:long_name = "day threshold compared against days since leaves became off-allometry" ;
	double fates_phen_drought_threshold ;
		fates_phen_drought_threshold:units = "m3/m3" ;
		fates_phen_drought_threshold:long_name = "liquid volume in soil layer, threashold for drought phenology" ;
	double fates_phen_mindayson ;
		fates_phen_mindayson:units = "days" ;
		fates_phen_mindayson:long_name = "day threshold compared against days since leaves became on-allometry" ;
	double fates_phen_ncolddayslim ;
		fates_phen_ncolddayslim:units = "days" ;
		fates_phen_ncolddayslim:long_name = "day threshold exceedance for temperature leaf-drop" ;
	double fates_q10_froz ;
		fates_q10_froz:units = "unitless" ;
		fates_q10_froz:long_name = "Q10 for frozen-soil respiration rates" ;
	double fates_q10_mr ;
		fates_q10_mr:units = "unitless" ;
		fates_q10_mr:long_name = "Q10 for maintenance respiration" ;
	double fates_soil_salinity ;
		fates_soil_salinity:units = "ppt" ;
		fates_soil_salinity:long_name = "soil salinity used for model when not coupled to dynamic soil salinity" ;

// global attributes:
		:history = "This file was made from FatesPFTIndexSwapper.py \n",
			" Input File = /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_temp0.nc \n",
			" Indices = [1, 1, 1]\n",
			" Wed Sep 08 2021, 11:21:28: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_pftname --val moist_trop_tree --PFT 1\n",
			" Wed Sep 08 2021, 11:21:28: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_pftname --val dry_trop_tree --PFT 2\n",
			" Wed Sep 08 2021, 11:21:29: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_pftname --val C4_Grass --PFT 3\n",
			" Wed Sep 08 2021, 11:21:29: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_allom_frbstor_repro --val 0.0 --allpfts\n",
			" Wed Sep 08 2021, 11:21:29: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_seed_suppl --val 0.0 --allpfts\n",
			" Wed Sep 08 2021, 11:21:29: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_branch_turnover --val 75\n",
			" Wed Sep 08 2021, 11:21:30: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_fire_alpha_SH --val 0.1487\n",
			" Wed Sep 08 2021, 11:21:30: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_fire_bark_scaler --val 0.0301\n",
			" Wed Sep 08 2021, 11:21:30: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_fire_crown_depth_frac --val 0.33\n",
			" Wed Sep 08 2021, 11:21:30: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_fire_crown_kill --val 1.0\n",
			" Wed Sep 08 2021, 11:21:31: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_grperc --val 0.30\n",
			" Wed Sep 08 2021, 11:21:31: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_leaf_long --val 1.4025\n",
			" Wed Sep 08 2021, 11:21:31: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_mort_hf_sm_threshold --val 0.025\n",
			" Wed Sep 08 2021, 11:21:31: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_seed_suppl --val 0.0\n",
			" Wed Sep 08 2021, 11:21:32: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_branch_turnover --val 75\n",
			" Wed Sep 08 2021, 11:21:32: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_fire_alpha_SH --val 0.06\n",
			" Wed Sep 08 2021, 11:21:32: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_fire_bark_scaler --val 0.1085\n",
			" Wed Sep 08 2021, 11:21:32: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_fire_crown_depth_frac --val 0.1\n",
			" Wed Sep 08 2021, 11:21:33: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_fire_crown_kill --val 0.05\n",
			" Wed Sep 08 2021, 11:21:33: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_grperc --val 0.30\n",
			" Wed Sep 08 2021, 11:21:33: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_leaf_long --val 1.4025\n",
			" Wed Sep 08 2021, 11:21:33: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_mort_hf_sm_threshold --val 0.025\n",
			" Wed Sep 08 2021, 11:21:34: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_seed_suppl --val 0.0\n",
			" Wed Sep 08 2021, 11:21:34: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_woody --val 0\n",
			" Wed Sep 08 2021, 11:21:34: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_alloc_storage_cushion --val 2.25\n",
			" Wed Sep 08 2021, 11:21:34: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_agb1 --val 0.000964\n",
			" Wed Sep 08 2021, 11:21:35: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_agb2 --val 1.9462\n",
			" Wed Sep 08 2021, 11:21:35: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_agb3 --val 0\n",
			" Wed Sep 08 2021, 11:21:35: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_agb4 --val 0\n",
			" Wed Sep 08 2021, 11:21:35: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_agb_frac --val 1\n",
			" Wed Sep 08 2021, 11:21:36: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_amode --val 1\n",
			" Wed Sep 08 2021, 11:21:36: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2bl1 --val 0.000964\n",
			" Wed Sep 08 2021, 11:21:36: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2bl2 --val 1.9492\n",
			" Wed Sep 08 2021, 11:21:36: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2bl3 --val 0\n",
			" Wed Sep 08 2021, 11:21:37: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2ca_coefficient_max --val 0.03\n",
			" Wed Sep 08 2021, 11:21:37: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2ca_coefficient_min --val 0.01\n",
			" Wed Sep 08 2021, 11:21:37: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2h1 --val 1\n",
			" Wed Sep 08 2021, 11:21:37: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2h2 --val 1\n",
			" Wed Sep 08 2021, 11:21:38: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_d2h3 --val -999.9\n",
			" Wed Sep 08 2021, 11:21:38: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_dbh_maxheight --val 1\n",
			" Wed Sep 08 2021, 11:21:38: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_hmode --val 3\n",
			" Wed Sep 08 2021, 11:21:38: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_la_per_sa_int --val 1000\n",
			" Wed Sep 08 2021, 11:21:39: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_l2fr --val 1\n",
			" Wed Sep 08 2021, 11:21:39: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_lmode --val 1\n",
			" Wed Sep 08 2021, 11:21:39: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_allom_sai_scaler --val 0.0012\n",
			" Wed Sep 08 2021, 11:21:40: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_branch_turnover --val 0.3208\n",
			" Wed Sep 08 2021, 11:21:40: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_fire_crown_depth_frac --val 1\n",
			" Wed Sep 08 2021, 11:21:40: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_fire_alpha_SH --val 1\n",
			" Wed Sep 08 2021, 11:21:40: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_fire_crown_kill --val 1\n",
			" Wed Sep 08 2021, 11:21:41: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_fnrt_prof_a --val 7\n",
			" Wed Sep 08 2021, 11:21:41: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_fnrt_prof_b --val 1\n",
			" Wed Sep 08 2021, 11:21:41: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_grperc --val 0.20\n",
			" Wed Sep 08 2021, 11:21:41: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_stomatal_slope_ballberry --val 4\n",
			" Wed Sep 08 2021, 11:21:42: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_clumping_index --val 0.85\n",
			" Wed Sep 08 2021, 11:21:42: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_c3psn --val 0\n",
			" Wed Sep 08 2021, 11:21:42: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_long --val 0.3208\n",
			" Wed Sep 08 2021, 11:21:42: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_stor_priority --val 0.8\n",
			" Wed Sep 08 2021, 11:21:43: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_slamax --val 0.02\n",
			" Wed Sep 08 2021, 11:21:43: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_slatop --val 0.02\n",
			" Wed Sep 08 2021, 11:21:43: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_xl --val -0.3\n",
			" Wed Sep 08 2021, 11:21:43: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_vcmax25top --val 30\n",
			" Wed Sep 08 2021, 11:21:44: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_prt_nitr_stoich_p1 --val .16,.024,1.e-8,1.e-8,0.,.0047\n",
			" Wed Sep 08 2021, 11:21:44: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_prt_phos_stoich_p1 --val .004,0024,1.e-9,1.e-9,0.,.00047\n",
			" Wed Sep 08 2021, 11:21:44: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_prt_phos_stoich_p2 --val .0033,0024,1.e-9,1.e-9,0.,.00047\n",
			" Wed Sep 08 2021, 11:21:44: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_mort_scalar_cstarvation --val 0.2\n",
			" Wed Sep 08 2021, 11:21:45: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_recruit_hgt_min --val 0.5\n",
			" Wed Sep 08 2021, 11:21:45: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_recruit_initd --val 20\n",
			" Wed Sep 08 2021, 11:21:45: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_seed_alloc --val 0.1\n",
			" Wed Sep 08 2021, 11:21:46: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_seed_alloc_mature --val 0.9\n",
			" Wed Sep 08 2021, 11:21:46: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_seed_dbh_repro_threshold --val 0.5\n",
			" Wed Sep 08 2021, 11:21:46: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_seed_suppl --val 0.0\n",
			" Wed Sep 08 2021, 11:21:46: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_wood_density --val 0.01\n",
			" Wed Sep 08 2021, 11:21:47: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rholnir --val 0.46 --PFT 1\n",
			" Wed Sep 08 2021, 11:21:47: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rholnir --val 0.46 --PFT 2\n",
			" Wed Sep 08 2021, 11:21:47: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rholnir --val 0.28 --PFT 3\n",
			" Wed Sep 08 2021, 11:21:48: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rholvis --val 0.11 --PFT 1\n",
			" Wed Sep 08 2021, 11:21:48: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rholvis --val 0.11 --PFT 2\n",
			" Wed Sep 08 2021, 11:21:49: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rholvis --val 0.05 --PFT 3\n",
			" Wed Sep 08 2021, 11:21:49: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rhosnir --val 0.49 --PFT 1\n",
			" Wed Sep 08 2021, 11:21:49: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rhosnir --val 0.49 --PFT 2\n",
			" Wed Sep 08 2021, 11:21:49: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rhosvis --val 0.21 --PFT 1\n",
			" Wed Sep 08 2021, 11:21:50: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_rhosvis --val 0.21 --PFT 2\n",
			" Wed Sep 08 2021, 11:21:50: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_taulnir --val 0.33 --PFT 1\n",
			" Wed Sep 08 2021, 11:21:50: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_taulnir --val 0.33 --PFT 2\n",
			" Wed Sep 08 2021, 11:21:50: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_taulnir --val 0.40 --PFT 3\n",
			" Wed Sep 08 2021, 11:21:51: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_taulvis --val 0.06 --PFT 1\n",
			" Wed Sep 08 2021, 11:21:51: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_taulvis --val 0.06 --PFT 2\n",
			" Wed Sep 08 2021, 11:21:51: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_taulvis --val 0.05 --PFT 3\n",
			" Wed Sep 08 2021, 11:21:51: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_fire_threshold --val 25\n",
			" Wed Sep 08 2021, 11:21:52: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_fire_drying_ratio --val 40000\n",
			" Wed Sep 08 2021, 11:21:52: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_history_sizeclass_bin_edges --val 0,5,10,15,20,30,40,50,60,70,80,90,100\n",
			" Wed Sep 08 2021, 11:21:52: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_wood_density --val 0.6305\n",
			" Wed Sep 08 2021, 11:21:52: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_wood_density --val 0.695\n",
			" Wed Sep 08 2021, 11:21:53: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_leaf_vcmax25top --val 41\n",
			" Wed Sep 08 2021, 11:21:53: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_leaf_vcmax25top --val 41\n",
			" Wed Sep 08 2021, 11:21:53: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 1 --var fates_prt_nitr_stoich_p1 --val .02674866,.024,1.e-8,1.e-8,0.,.0047\n",
			" Wed Sep 08 2021, 11:21:53: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 2 --var fates_prt_nitr_stoich_p1 --val .02674866,.024,1.e-8,1.e-8,0.,.0047\n",
			" Wed Sep 08 2021, 11:21:54: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_vcmax25top --val 40\n",
			" Wed Sep 08 2021, 11:21:54: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_grperc --val 0.11\n",
			" Wed Sep 08 2021, 11:21:54: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_slamax --val 0.0135\n",
			" Wed Sep 08 2021, 11:21:54: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_leaf_slatop --val 0.0135\n",
			" Wed Sep 08 2021, 11:21:55: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --PFT 3 --var fates_prt_nitr_stoich_p1 --val .16,.024,1.e-8,1.e-8,0.,.0047\n",
			" Wed Sep 08 2021, 11:21:55: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_fire_FBD --val 15.4,16.8,19.6,999,4,0.95\n",
			" Wed Sep 08 2021, 11:21:55: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_fire_drying_ratio --val 66000\n",
			" Wed Sep 08 2021, 11:21:55: modify_fates_paramfile.py --O --fin /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --fout /glade/work/jkshuman/FATES_data/parameter_files/C4Gr_TropTrees/param_file_cg_BDliveG1_66dry_C4sla0135_nitr16C4_grresp11_vcmx40_wooddens_fireparams_nitr_BCIens_vcmxtrees41_C440_storcush12_leaflong_grwresp30_75branch_25thresh_20210908.nc --var fates_fire_cg_strikes --val 0.1" ;
data:

 fates_history_sizeclass_bin_edges = 0, 5, 10, 15, 20, 30, 40, 50, 60, 70, 
    80, 90, 100 ;

 fates_history_ageclass_bin_edges = 0, 1, 2, 5, 10, 20, 50 ;

 fates_prt_organ_name =
  "leaf                                             ",
  "fine root                                        ",
  "sapwood                                          ",
  "storage                                          ",
  "reproduction                                     ",
  "structure                                        " ;

 fates_prt_alloc_priority =
  1, 1, 1,
  2, 2, 2,
  3, 3, 3,
  3, 3, 3,
  0, 0, 0,
  4, 4, 4 ;

 fates_prt_nitr_stoich_p1 =
  0.0267486590892076, 0.0267486590892076, 0.159999996423721,
  0.0240000002086163, 0.0240000002086163, 0.0240000002086163,
  9.99999993922529e-09, 9.99999993922529e-09, 9.99999993922529e-09,
  9.99999993922529e-09, 9.99999993922529e-09, 9.99999993922529e-09,
  0, 0, 0,
  0.00469999993219972, 0.00469999993219972, 0.00469999993219972 ;

 fates_prt_nitr_stoich_p2 =
  0.033, 0.033, 0.033,
  0.024, 0.024, 0.024,
  1e-08, 1e-08, 1e-08,
  1e-08, 1e-08, 1e-08,
  0, 0, 0,
  0.0047, 0.0047, 0.0047 ;

 fates_prt_phos_stoich_p1 =
  0.0033, 0.0033, 0.00400000018998981,
  0.0024, 0.0024, 24,
  1e-09, 1e-09, 9.99999971718069e-10,
  1e-09, 1e-09, 9.99999971718069e-10,
  0, 0, 0,
  0.00047, 0.00047, 0.000469999999040738 ;

 fates_prt_phos_stoich_p2 =
  0.0033, 0.0033, 0.00329999998211861,
  0.0024, 0.0024, 24,
  1e-09, 1e-09, 9.99999971718069e-10,
  1e-09, 1e-09, 9.99999971718069e-10,
  0, 0, 0,
  0.00047, 0.00047, 0.000469999999040738 ;

 fates_turnover_carb_retrans =
  0.025, 0.025, 0.025,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0 ;

 fates_turnover_nitr_retrans =
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _ ;

 fates_turnover_phos_retrans =
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _ ;

 fates_fire_FBD = 15.3999996185303, 16.7999992370605, 19.6000003814697, 999, 
    4, 0.949999988079071 ;

 fates_fire_SAV = 13, 3.58, 0.98, 0.2, 66, 66 ;

 fates_fire_low_moisture_Coeff = 1.12, 1.09, 0.98, 0.8, 1.15, 1.15 ;

 fates_fire_low_moisture_Slope = 0.62, 0.72, 0.85, 0.8, 0.62, 0.62 ;

 fates_fire_mid_moisture = 0.72, 0.51, 0.38, 1, 0.8, 0.8 ;

 fates_fire_mid_moisture_Coeff = 2.35, 1.47, 1.06, 0.8, 3.2, 3.2 ;

 fates_fire_mid_moisture_Slope = 2.35, 1.47, 1.06, 0.8, 3.2, 3.2 ;

 fates_fire_min_moisture = 0.18, 0.12, 0, 0, 0.24, 0.24 ;

 fates_history_height_bin_edges = 0, 0.1, 0.3, 1, 3, 10 ;

 fates_max_decomp = 0.52, 0.383, 0.383, 0.19, 1, 999 ;

 fates_hydr_avuln_node =
  2, 2, 2,
  2, 2, 2,
  2, 2, 2,
  2, 2, 2 ;

 fates_hydr_epsil_node =
  12, 12, 12,
  10, 10, 10,
  10, 10, 10,
  8, 8, 8 ;

 fates_hydr_fcap_node =
  0, 0, 0,
  0.08, 0.08, 0.08,
  0.08, 0.08, 0.08,
  0, 0, 0 ;

 fates_hydr_kmax_node =
  -999, -999, -999,
  3, 3, 3,
  -999, -999, -999,
  -999, -999, -999 ;

 fates_hydr_p50_node =
  -2.25, -2.25, -2.25,
  -2.25, -2.25, -2.25,
  -2.25, -2.25, -2.25,
  -2.25, -2.25, -2.25 ;

 fates_hydr_pinot_node =
  -1.465984, -1.465984, -1.465984,
  -1.22807, -1.22807, -1.22807,
  -1.22807, -1.22807, -1.22807,
  -1.043478, -1.043478, -1.043478 ;

 fates_hydr_pitlp_node =
  -1.67, -1.67, -1.67,
  -1.4, -1.4, -1.4,
  -1.4, -1.4, -1.4,
  -1.2, -1.2, -1.2 ;

 fates_hydr_resid_node =
  0.16, 0.16, 0.16,
  0.21, 0.21, 0.21,
  0.21, 0.21, 0.21,
  0.11, 0.11, 0.11 ;

 fates_hydr_thetas_node =
  0.65, 0.65, 0.65,
  0.65, 0.65, 0.65,
  0.65, 0.65, 0.65,
  0.75, 0.75, 0.75 ;

 fates_CWD_frac = 0.045, 0.075, 0.21, 0.67 ;

 fates_pftname =
  "moist_trop_tree                                             ",
  "dry_trop_tree                                               ",
  "C4_Grass                                                    " ;

 fates_alloc_storage_cushion = 1.2, 1.2, 2.25 ;

 fates_allom_agb1 = 0.0673, 0.0673, 0.000964 ;

 fates_allom_agb2 = 0.976, 0.976, 1.9462 ;

 fates_allom_agb3 = _, _, 0 ;

 fates_allom_agb4 = _, _, 0 ;

 fates_allom_agb_frac = 0.6, 0.6, 1 ;

 fates_allom_amode = 3, 3, 1 ;

 fates_allom_blca_expnt_diff = 0, 0, 0 ;

 fates_allom_cmode = 1, 1, 1 ;

 fates_allom_d2bl1 = 0.1266844, 0.1266844, 0.000964 ;

 fates_allom_d2bl2 = 1.281329, 1.281329, 1.9492 ;

 fates_allom_d2bl3 = _, _, 0 ;

 fates_allom_d2ca_coefficient_max = 0.768654, 0.768654, 0.03 ;

 fates_allom_d2ca_coefficient_min = 0.768654, 0.768654, 0.01 ;

 fates_allom_d2h1 = 57.6, 57.6, 1 ;

 fates_allom_d2h2 = 0.74, 0.74, 1 ;

 fates_allom_d2h3 = 21.6, 21.6, -999.9 ;

 fates_allom_dbh_maxheight = 200, 200, 1 ;

 fates_allom_fmode = 2, 2, 2 ;

 fates_allom_frbstor_repro = 0, 0, 0 ;

 fates_allom_hmode = 5, 5, 3 ;

 fates_allom_l2fr = 0.4863088, 0.4863088, 1 ;

 fates_allom_la_per_sa_int = 0.8, 0.8, 1000 ;

 fates_allom_la_per_sa_slp = 0, 0, 0 ;

 fates_allom_lmode = 3, 3, 1 ;

 fates_allom_sai_scaler = 0.1, 0.1, 0.0012 ;

 fates_allom_smode = 1, 1, 1 ;

 fates_allom_stmode = 1, 1, 1 ;

 fates_branch_turnover = 75, 75, 0.3208 ;

 fates_c2b = 2, 2, 2 ;

 fates_displar = 0.67, 0.67, 0.67 ;

 fates_eca_alpha_ptase = 0.5, 0.5, 0.5 ;

 fates_eca_decompmicc = 280, 280, 280 ;

 fates_eca_km_nh4 = 0.14, 0.14, 0.14 ;

 fates_eca_km_no3 = 0.27, 0.27, 0.27 ;

 fates_eca_km_p = 0.1, 0.1, 0.1 ;

 fates_eca_km_ptase = 1, 1, 1 ;

 fates_eca_lambda_ptase = 1, 1, 1 ;

 fates_eca_vmax_nh4 = 1.5e-07, 1.5e-07, 1.5e-07 ;

 fates_eca_vmax_no3 = 1.5e-08, 1.5e-08, 1.5e-08 ;

 fates_eca_vmax_p = 1.5e-09, 1.5e-09, 1.5e-09 ;

 fates_eca_vmax_ptase = 5e-09, 5e-09, 5e-09 ;

 fates_fire_alpha_SH = 0.1487, 0.06, 1 ;

 fates_fire_bark_scaler = 0.0301, 0.1085, 0.07 ;

 fates_fire_crown_depth_frac = 0.33, 0.1, 1 ;

 fates_fire_crown_kill = 1, 0.05, 1 ;

 fates_fnrt_prof_a = 7, 7, 7 ;

 fates_fnrt_prof_b = 1, 1, 1 ;

 fates_fnrt_prof_mode = 3, 3, 3 ;

 fates_fr_fcel = 0.5, 0.5, 0.5 ;

 fates_fr_flab = 0.25, 0.25, 0.25 ;

 fates_fr_flig = 0.25, 0.25, 0.25 ;

 fates_grperc = 0.3, 0.3, 0.11 ;

 fates_hydr_avuln_gs = 2.5, 2.5, 2.5 ;

 fates_hydr_p50_gs = -1.5, -1.5, -1.5 ;

 fates_hydr_p_taper = 0.333, 0.333, 0.333 ;

 fates_hydr_rfrac_stem = 0.625, 0.625, 0.625 ;

 fates_hydr_rs2 = 0.0001, 0.0001, 0.0001 ;

 fates_hydr_srl = 25, 25, 25 ;

 fates_leaf_c3psn = 1, 1, 0 ;

 fates_leaf_clumping_index = 0.85, 0.85, 0.85 ;

 fates_leaf_diameter = 0.04, 0.04, 0.04 ;

 fates_leaf_jmaxha = 43540, 43540, 43540 ;

 fates_leaf_jmaxhd = 152040, 152040, 152040 ;

 fates_leaf_jmaxse = 495, 495, 495 ;

 fates_leaf_slamax = 0.03991654, 0.03991654, 0.0135 ;

 fates_leaf_slatop = 0.01995827, 0.01995827, 0.0135 ;

 fates_leaf_stomatal_intercept = 10000, 10000, 10000 ;

 fates_leaf_stomatal_slope_ballberry = 8, 8, 4 ;

 fates_leaf_stomatal_slope_medlyn = 4.1, 4.1, 4.1 ;

 fates_leaf_stor_priority = 0.8, 0.8, 0.8 ;

 fates_leaf_tpuha = 53100, 53100, 53100 ;

 fates_leaf_tpuhd = 150650, 150650, 150650 ;

 fates_leaf_tpuse = 490, 490, 490 ;

 fates_leaf_vcmaxha = 65330, 65330, 65330 ;

 fates_leaf_vcmaxhd = 149250, 149250, 149250 ;

 fates_leaf_vcmaxse = 485, 485, 485 ;

 fates_leaf_xl = 0.1, 0.1, -0.3 ;

 fates_lf_fcel = 0.5, 0.5, 0.5 ;

 fates_lf_flab = 0.25, 0.25, 0.25 ;

 fates_lf_flig = 0.25, 0.25, 0.25 ;

 fates_maintresp_reduction_curvature = 0.01, 0.01, 0.01 ;

 fates_maintresp_reduction_intercept = 1, 1, 1 ;

 fates_mort_bmort = 0.01303514, 0.01303514, 0.01303514 ;

 fates_mort_freezetol = 2.5, 2.5, 2.5 ;

 fates_mort_hf_flc_threshold = 0.5, 0.5, 0.5 ;

 fates_mort_hf_sm_threshold = 0.025, 0.025, 1e-06 ;

 fates_mort_ip_age_senescence = _, _, _ ;

 fates_mort_ip_size_senescence = _, _, _ ;

 fates_mort_r_age_senescence = _, _, _ ;

 fates_mort_r_size_senescence = _, _, _ ;

 fates_mort_scalar_coldstress = 3, 3, 3 ;

 fates_mort_scalar_cstarvation = 0.02955703, 0.02955703, 0.2 ;

 fates_mort_scalar_hydrfailure = 0.6, 0.6, 0.6 ;

 fates_nfix1 = _, _, _ ;

 fates_nfix2 = _, _, _ ;

 fates_phen_cold_size_threshold = 0, 0, 0 ;

 fates_phen_evergreen = 1, 1, 1 ;

 fates_phen_season_decid = 0, 0, 0 ;

 fates_phen_stem_drop_fraction = 0, 0, 0 ;

 fates_phen_stress_decid = 0, 0, 0 ;

 fates_phenflush_fraction = _, _, _ ;

 fates_prescribed_mortality_canopy = 0.0194, 0.0194, 0.0194 ;

 fates_prescribed_mortality_understory = 0.025, 0.025, 0.025 ;

 fates_prescribed_npp_canopy = 0.4, 0.4, 0.4 ;

 fates_prescribed_npp_understory = 0.03125, 0.03125, 0.03125 ;

 fates_prescribed_nuptake = 5, 5, 5 ;

 fates_prescribed_puptake = 5, 5, 5 ;

 fates_prescribed_recruitment = 0.02, 0.02, 0.02 ;

 fates_recruit_hgt_min = 1.3, 1.3, 0.5 ;

 fates_recruit_initd = 0.2, 0.2, 20 ;

 fates_rholnir = 0.46, 0.46, 0.28 ;

 fates_rholvis = 0.11, 0.11, 0.05 ;

 fates_rhosnir = 0.49, 0.49, 0.39 ;

 fates_rhosvis = 0.21, 0.21, 0.16 ;

 fates_root_long = 1, 1, 1 ;

 fates_seed_alloc = 0.04680188, 0.04680188, 0.1 ;

 fates_seed_alloc_mature = 0, 0, 0.9 ;

 fates_seed_dbh_repro_threshold = 150, 150, 0.5 ;

 fates_seed_decay_rate = 0.51, 0.51, 0.51 ;

 fates_seed_germination_rate = 0.5, 0.5, 0.5 ;

 fates_seed_suppl = 0, 0, 0 ;

 fates_senleaf_long_fdrought = 1, 1, 1 ;

 fates_smpsc = -255000, -255000, -255000 ;

 fates_smpso = -66000, -66000, -66000 ;

 fates_taulnir = 0.33, 0.33, 0.4 ;

 fates_taulvis = 0.06, 0.06, 0.05 ;

 fates_tausnir = 0.001, 0.001, 0.001 ;

 fates_tausvis = 0.001, 0.001, 0.001 ;

 fates_trim_inc = 0.03, 0.03, 0.03 ;

 fates_trim_limit = 0.3, 0.3, 0.3 ;

 fates_turnover_retrans_mode = 1, 1, 1 ;

 fates_wood_density = 0.6305, 0.695, 0.01 ;

 fates_woody = 1, 1, 0 ;

 fates_z0mr = 0.055, 0.055, 0.055 ;

 fates_history_coageclass_bin_edges = 0, 5 ;

 fates_leaf_long =
  1.4025, 1.4025, 0.3208 ;

 fates_leaf_vcmax25top =
  41, 41, 40 ;

 fates_base_mr_20 = 2.52e-06 ;

 fates_canopy_closure_thresh = 0.8 ;

 fates_cohort_age_fusion_tol = 0.08 ;

 fates_cohort_size_fusion_tol = 0.08 ;

 fates_comp_excln = -1 ;

 fates_cwd_fcel = 0.76 ;

 fates_cwd_flig = 0.24 ;

 fates_eca_plant_escalar = 1.25e-05 ;

 fates_fire_active_crown_fire = 0 ;

 fates_fire_cg_strikes = 0.1 ;

 fates_fire_drying_ratio = 66000 ;

 fates_fire_durat_slope = -11.06 ;

 fates_fire_fdi_a = 17.62 ;

 fates_fire_fdi_alpha = 0.00037 ;

 fates_fire_fdi_b = 243.12 ;

 fates_fire_fuel_energy = 18000 ;

 fates_fire_max_durat = 240 ;

 fates_fire_miner_damp = 0.41739 ;

 fates_fire_miner_total = 0.055 ;

 fates_fire_nignitions = 15 ;

 fates_fire_part_dens = 513 ;

 fates_fire_threshold = 25 ;

 fates_hydr_kmax_rsurf1 = 20 ;

 fates_hydr_kmax_rsurf2 = 0.0001 ;

 fates_hydr_psi0 = 0 ;

 fates_hydr_psicap = -0.6 ;

 fates_init_litter = 0.05 ;

 fates_leaf_stomatal_model = 1 ;

 fates_logging_coll_under_frac = 0.55983 ;

 fates_logging_collateral_frac = 0.05 ;

 fates_logging_dbhmax = _ ;

 fates_logging_dbhmax_infra = 35 ;

 fates_logging_dbhmin = 50 ;

 fates_logging_direct_frac = 0.15 ;

 fates_logging_event_code = -30 ;

 fates_logging_export_frac = 0.8 ;

 fates_logging_mechanical_frac = 0.05 ;

 fates_mort_disturb_frac = 0.5 ;

 fates_mort_understorey_death = 1 ;

 fates_patch_fusion_tol = 0.05 ;

 fates_phen_a = -68 ;

 fates_phen_b = 638 ;

 fates_phen_c = -0.01 ;

 fates_phen_chiltemp = 5 ;

 fates_phen_coldtemp = 7.5 ;

 fates_phen_doff_time = 100 ;

 fates_phen_drought_threshold = 0.15 ;

 fates_phen_mindayson = 90 ;

 fates_phen_ncolddayslim = 5 ;

 fates_q10_froz = 1.5 ;

 fates_q10_mr = 1.5 ;

 fates_soil_salinity = 0.4 ;
}
